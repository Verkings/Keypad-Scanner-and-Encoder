
module fifo_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;
  wire   [31:2] carry;

  CHA1X1 U1_1_30 ( .A(A[30]), .B(n23), .CO(carry[31]), .S(SUM[30]) );
  CHA1X1 U1_1_16 ( .A(A[16]), .B(n1), .CO(carry[17]), .S(SUM[16]) );
  CHA1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CHA1X2 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  CHA1X2 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  CHA1X2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CHA1X2 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  CHA1X2 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  CHA1X2 U1_1_12 ( .A(A[12]), .B(n11), .CO(carry[13]), .S(SUM[12]) );
  CIVX1 U1 ( .A(n39), .Z(carry[15]) );
  CNR2IX2 U2 ( .B(A[15]), .A(n39), .Z(n1) );
  CND2IX2 U3 ( .B(n2), .A(carry[13]), .Z(n6) );
  CIVX20 U4 ( .A(A[13]), .Z(n2) );
  CIVXL U5 ( .A(n41), .Z(carry[21]) );
  CIVX2 U6 ( .A(n6), .Z(n3) );
  CIVXL U7 ( .A(n6), .Z(carry[14]) );
  CIVX2 U8 ( .A(n18), .Z(n4) );
  CIVXL U9 ( .A(n18), .Z(carry[19]) );
  CEOXL U10 ( .A(A[19]), .B(carry[19]), .Z(SUM[19]) );
  CIVX4 U11 ( .A(n5), .Z(carry[20]) );
  CND2X2 U12 ( .A(n4), .B(A[19]), .Z(n5) );
  CEOXL U13 ( .A(A[13]), .B(carry[13]), .Z(SUM[13]) );
  CEOXL U14 ( .A(A[15]), .B(carry[15]), .Z(SUM[15]) );
  CND2IX4 U15 ( .B(n40), .A(carry[20]), .Z(n41) );
  CNR2IX4 U16 ( .B(A[27]), .A(n20), .Z(n8) );
  CND2IX2 U17 ( .B(n7), .A(carry[26]), .Z(n20) );
  CIVX20 U18 ( .A(A[26]), .Z(n7) );
  CIVX2 U19 ( .A(n42), .Z(n9) );
  CIVXL U20 ( .A(n42), .Z(n33) );
  CNR2IX4 U21 ( .B(A[21]), .A(n41), .Z(n10) );
  CNR2IX2 U22 ( .B(A[11]), .A(n17), .Z(n11) );
  CEOXL U23 ( .A(A[2]), .B(n33), .Z(SUM[2]) );
  CND2X2 U24 ( .A(n9), .B(A[2]), .Z(n12) );
  CIVX2 U25 ( .A(n12), .Z(carry[3]) );
  CND2X2 U26 ( .A(carry[3]), .B(A[3]), .Z(n43) );
  CIVXL U27 ( .A(n20), .Z(carry[27]) );
  CIVXL U28 ( .A(n17), .Z(carry[11]) );
  CND2IX2 U29 ( .B(n13), .A(carry[18]), .Z(n18) );
  CIVX20 U30 ( .A(A[18]), .Z(n13) );
  CIVXL U31 ( .A(n33), .Z(n14) );
  CIVXL U32 ( .A(carry[21]), .Z(n15) );
  CIVX2 U33 ( .A(n15), .Z(n16) );
  CEOXL U34 ( .A(A[10]), .B(carry[10]), .Z(SUM[10]) );
  CND2X2 U35 ( .A(A[10]), .B(carry[10]), .Z(n17) );
  CEOXL U36 ( .A(A[18]), .B(carry[18]), .Z(SUM[18]) );
  CEOXL U37 ( .A(A[5]), .B(carry[5]), .Z(SUM[5]) );
  CIVX2 U38 ( .A(n19), .Z(carry[6]) );
  CND2X2 U39 ( .A(A[5]), .B(carry[5]), .Z(n19) );
  CEOXL U40 ( .A(A[26]), .B(carry[26]), .Z(SUM[26]) );
  CIVX1 U41 ( .A(n25), .Z(carry[29]) );
  CND2IX2 U42 ( .B(n21), .A(carry[8]), .Z(n27) );
  CIVX20 U43 ( .A(A[8]), .Z(n21) );
  CND2IX2 U44 ( .B(n22), .A(n35), .Z(n26) );
  CIVX20 U45 ( .A(A[24]), .Z(n22) );
  CNR2IX2 U46 ( .B(A[29]), .A(n25), .Z(n23) );
  CDLY1XL U47 ( .A(n14), .Z(n24) );
  CEOXL U48 ( .A(A[28]), .B(n8), .Z(SUM[28]) );
  CND2X2 U49 ( .A(n8), .B(A[28]), .Z(n25) );
  CEOXL U50 ( .A(A[24]), .B(n35), .Z(SUM[24]) );
  CIVX2 U51 ( .A(n26), .Z(carry[25]) );
  CEOXL U52 ( .A(A[8]), .B(carry[8]), .Z(SUM[8]) );
  CIVX2 U53 ( .A(n27), .Z(carry[9]) );
  CEOXL U54 ( .A(A[21]), .B(n16), .Z(SUM[21]) );
  CNR2X4 U55 ( .A(n37), .B(n36), .Z(n35) );
  CND2X4 U56 ( .A(A[22]), .B(n10), .Z(n37) );
  CND2X1 U57 ( .A(carry[31]), .B(n32), .Z(n30) );
  CND2X2 U58 ( .A(n28), .B(n29), .Z(n31) );
  CND2X2 U59 ( .A(n31), .B(n30), .Z(SUM[31]) );
  CIVX1 U60 ( .A(carry[31]), .Z(n28) );
  CIVX2 U61 ( .A(n32), .Z(n29) );
  CIVXL U62 ( .A(A[31]), .Z(n32) );
  CIVXL U63 ( .A(A[0]), .Z(SUM[0]) );
  CIVXL U64 ( .A(n24), .Z(carry[2]) );
  CND2IX2 U65 ( .B(n34), .A(n3), .Z(n39) );
  CIVX20 U66 ( .A(A[14]), .Z(n34) );
  CIVX20 U67 ( .A(A[23]), .Z(n36) );
  CEOXL U68 ( .A(A[22]), .B(n10), .Z(SUM[22]) );
  CIVX3 U69 ( .A(n37), .Z(carry[23]) );
  CEOXL U70 ( .A(A[23]), .B(carry[23]), .Z(SUM[23]) );
  CEOXL U71 ( .A(A[29]), .B(carry[29]), .Z(SUM[29]) );
  CEOXL U72 ( .A(A[11]), .B(carry[11]), .Z(SUM[11]) );
  CAN2XL U73 ( .A(A[2]), .B(carry[2]), .Z(n38) );
  CEOXL U74 ( .A(A[14]), .B(carry[14]), .Z(SUM[14]) );
  CIVX20 U75 ( .A(A[20]), .Z(n40) );
  CEOXL U76 ( .A(A[20]), .B(carry[20]), .Z(SUM[20]) );
  CEOXL U77 ( .A(A[1]), .B(A[0]), .Z(SUM[1]) );
  CND2X2 U78 ( .A(A[1]), .B(A[0]), .Z(n42) );
  CEOXL U79 ( .A(A[3]), .B(n38), .Z(SUM[3]) );
  CIVX2 U80 ( .A(n43), .Z(carry[4]) );
  CEOXL U81 ( .A(A[27]), .B(carry[27]), .Z(SUM[27]) );
endmodule


module fifo_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B_not[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [32:0] carry;

  CENX1 U1 ( .A(A[30]), .B(carry[30]), .Z(DIFF[30]) );
  CND2IX2 U2 ( .B(\B_not[0] ), .A(n55), .Z(carry[1]) );
  CND2IX2 U3 ( .B(A[10]), .A(n1), .Z(carry[11]) );
  CND2IX2 U4 ( .B(A[11]), .A(n2), .Z(carry[12]) );
  CND2IX2 U5 ( .B(A[16]), .A(n11), .Z(carry[17]) );
  CND2IX2 U6 ( .B(A[18]), .A(n14), .Z(carry[19]) );
  CND2IX2 U7 ( .B(A[23]), .A(n25), .Z(carry[24]) );
  CND2IX2 U8 ( .B(A[24]), .A(n26), .Z(carry[25]) );
  CENXL U9 ( .A(A[26]), .B(carry[26]), .Z(DIFF[26]) );
  CENXL U10 ( .A(A[3]), .B(carry[3]), .Z(DIFF[3]) );
  CENXL U11 ( .A(A[17]), .B(carry[17]), .Z(DIFF[17]) );
  CENXL U12 ( .A(A[12]), .B(carry[12]), .Z(DIFF[12]) );
  CENXL U13 ( .A(A[7]), .B(carry[7]), .Z(DIFF[7]) );
  CENXL U14 ( .A(A[4]), .B(carry[4]), .Z(DIFF[4]) );
  CENXL U15 ( .A(A[5]), .B(carry[5]), .Z(DIFF[5]) );
  CENXL U16 ( .A(A[19]), .B(carry[19]), .Z(DIFF[19]) );
  CENXL U17 ( .A(A[18]), .B(carry[18]), .Z(DIFF[18]) );
  CENXL U18 ( .A(A[25]), .B(carry[25]), .Z(DIFF[25]) );
  CENXL U19 ( .A(A[13]), .B(carry[13]), .Z(DIFF[13]) );
  CENXL U20 ( .A(A[14]), .B(carry[14]), .Z(DIFF[14]) );
  CENXL U21 ( .A(A[9]), .B(carry[9]), .Z(DIFF[9]) );
  CENXL U22 ( .A(A[8]), .B(carry[8]), .Z(DIFF[8]) );
  CENXL U23 ( .A(A[2]), .B(carry[2]), .Z(DIFF[2]) );
  CENXL U24 ( .A(A[21]), .B(carry[21]), .Z(DIFF[21]) );
  CENXL U25 ( .A(A[28]), .B(carry[28]), .Z(DIFF[28]) );
  CENXL U26 ( .A(A[20]), .B(carry[20]), .Z(DIFF[20]) );
  CENXL U27 ( .A(A[16]), .B(carry[16]), .Z(DIFF[16]) );
  CENXL U28 ( .A(A[27]), .B(carry[27]), .Z(DIFF[27]) );
  CENXL U29 ( .A(A[15]), .B(carry[15]), .Z(DIFF[15]) );
  CENXL U30 ( .A(A[10]), .B(carry[10]), .Z(DIFF[10]) );
  CENXL U31 ( .A(A[11]), .B(carry[11]), .Z(DIFF[11]) );
  CENXL U32 ( .A(\B_not[0] ), .B(A[0]), .Z(DIFF[0]) );
  CENXL U33 ( .A(A[1]), .B(carry[1]), .Z(DIFF[1]) );
  CIVXL U34 ( .A(A[29]), .Z(n35) );
  CENXL U35 ( .A(A[23]), .B(carry[23]), .Z(DIFF[23]) );
  CENXL U36 ( .A(A[24]), .B(carry[24]), .Z(DIFF[24]) );
  CENXL U37 ( .A(A[29]), .B(carry[29]), .Z(DIFF[29]) );
  CENXL U38 ( .A(A[6]), .B(carry[6]), .Z(DIFF[6]) );
  CIVXL U39 ( .A(A[22]), .Z(n23) );
  CENXL U40 ( .A(A[22]), .B(carry[22]), .Z(DIFF[22]) );
  CIVXL U41 ( .A(A[30]), .Z(n39) );
  CENXL U42 ( .A(A[31]), .B(carry[31]), .Z(DIFF[31]) );
  CIVX2 U43 ( .A(carry[10]), .Z(n1) );
  CIVX2 U44 ( .A(carry[11]), .Z(n2) );
  CND2X2 U45 ( .A(n3), .B(n4), .Z(carry[13]) );
  CIVX2 U46 ( .A(A[12]), .Z(n3) );
  CIVX2 U47 ( .A(carry[12]), .Z(n4) );
  CND2X2 U48 ( .A(n5), .B(n6), .Z(carry[14]) );
  CIVX2 U49 ( .A(A[13]), .Z(n5) );
  CIVX2 U50 ( .A(carry[13]), .Z(n6) );
  CND2X2 U51 ( .A(n7), .B(n8), .Z(carry[15]) );
  CIVX2 U52 ( .A(A[14]), .Z(n7) );
  CIVX2 U53 ( .A(carry[14]), .Z(n8) );
  CND2X2 U54 ( .A(n9), .B(n10), .Z(carry[16]) );
  CIVX2 U55 ( .A(A[15]), .Z(n9) );
  CIVX2 U56 ( .A(carry[15]), .Z(n10) );
  CIVX2 U57 ( .A(carry[16]), .Z(n11) );
  CND2X2 U58 ( .A(n12), .B(n13), .Z(carry[18]) );
  CIVX2 U59 ( .A(A[17]), .Z(n12) );
  CIVX2 U60 ( .A(carry[17]), .Z(n13) );
  CIVX2 U61 ( .A(carry[18]), .Z(n14) );
  CND2X2 U62 ( .A(n15), .B(n16), .Z(carry[20]) );
  CIVX2 U63 ( .A(A[19]), .Z(n15) );
  CIVX2 U64 ( .A(carry[19]), .Z(n16) );
  CND2X2 U65 ( .A(n17), .B(n18), .Z(carry[2]) );
  CIVX2 U66 ( .A(A[1]), .Z(n17) );
  CIVX2 U67 ( .A(carry[1]), .Z(n18) );
  CND2X2 U68 ( .A(n19), .B(n20), .Z(carry[21]) );
  CIVX2 U69 ( .A(A[20]), .Z(n19) );
  CIVX2 U70 ( .A(carry[20]), .Z(n20) );
  CND2X2 U71 ( .A(n21), .B(n22), .Z(carry[22]) );
  CIVX2 U72 ( .A(A[21]), .Z(n21) );
  CIVX2 U73 ( .A(carry[21]), .Z(n22) );
  CND2X2 U74 ( .A(n23), .B(n24), .Z(carry[23]) );
  CIVX2 U75 ( .A(carry[22]), .Z(n24) );
  CIVX2 U76 ( .A(carry[23]), .Z(n25) );
  CIVX2 U77 ( .A(carry[24]), .Z(n26) );
  CND2X2 U78 ( .A(n27), .B(n28), .Z(carry[26]) );
  CIVX2 U79 ( .A(A[25]), .Z(n27) );
  CIVX2 U80 ( .A(carry[25]), .Z(n28) );
  CND2X2 U81 ( .A(n29), .B(n30), .Z(carry[27]) );
  CIVX2 U82 ( .A(A[26]), .Z(n29) );
  CIVX2 U83 ( .A(carry[26]), .Z(n30) );
  CND2X2 U84 ( .A(n31), .B(n32), .Z(carry[28]) );
  CIVX2 U85 ( .A(A[27]), .Z(n31) );
  CIVX2 U86 ( .A(carry[27]), .Z(n32) );
  CND2X2 U87 ( .A(n33), .B(n34), .Z(carry[29]) );
  CIVX2 U88 ( .A(A[28]), .Z(n33) );
  CIVX2 U89 ( .A(carry[28]), .Z(n34) );
  CND2X2 U90 ( .A(n35), .B(n36), .Z(carry[30]) );
  CIVX2 U91 ( .A(carry[29]), .Z(n36) );
  CND2X2 U92 ( .A(n37), .B(n38), .Z(carry[3]) );
  CIVX2 U93 ( .A(A[2]), .Z(n37) );
  CIVX2 U94 ( .A(carry[2]), .Z(n38) );
  CND2X2 U95 ( .A(n39), .B(n40), .Z(carry[31]) );
  CIVX2 U96 ( .A(carry[30]), .Z(n40) );
  CND2X2 U97 ( .A(n41), .B(n42), .Z(carry[4]) );
  CIVX2 U98 ( .A(A[3]), .Z(n41) );
  CIVX2 U99 ( .A(carry[3]), .Z(n42) );
  CND2X2 U100 ( .A(n43), .B(n44), .Z(carry[5]) );
  CIVX2 U101 ( .A(A[4]), .Z(n43) );
  CIVX2 U102 ( .A(carry[4]), .Z(n44) );
  CND2X2 U103 ( .A(n45), .B(n46), .Z(carry[6]) );
  CIVX2 U104 ( .A(A[5]), .Z(n45) );
  CIVX2 U105 ( .A(carry[5]), .Z(n46) );
  CND2X2 U106 ( .A(n47), .B(n48), .Z(carry[7]) );
  CIVX2 U107 ( .A(A[6]), .Z(n47) );
  CIVX2 U108 ( .A(carry[6]), .Z(n48) );
  CND2X2 U109 ( .A(n49), .B(n50), .Z(carry[8]) );
  CIVX2 U110 ( .A(A[7]), .Z(n49) );
  CIVX2 U111 ( .A(carry[7]), .Z(n50) );
  CND2X2 U112 ( .A(n51), .B(n52), .Z(carry[9]) );
  CIVX2 U113 ( .A(A[8]), .Z(n51) );
  CIVX2 U114 ( .A(carry[8]), .Z(n52) );
  CND2X2 U115 ( .A(n53), .B(n54), .Z(carry[10]) );
  CIVX2 U116 ( .A(A[9]), .Z(n53) );
  CIVX2 U117 ( .A(carry[9]), .Z(n54) );
  CIVX2 U118 ( .A(A[0]), .Z(n55) );
  CIVX1 U119 ( .A(B[0]), .Z(\B_not[0] ) );
endmodule


module fifo ( code, full, empty, data, rd_enable, wr_enable, reset, clock );
  output [3:0] code;
  input [3:0] data;
  input rd_enable, wr_enable, reset, clock;
  output full, empty;
  wire   N1, N3, N4, N6, N7, N51, \memory[31][3] , \memory[31][2] ,
         \memory[31][1] , \memory[31][0] , \memory[30][3] , \memory[30][2] ,
         \memory[30][1] , \memory[30][0] , \memory[29][3] , \memory[29][2] ,
         \memory[29][1] , \memory[29][0] , \memory[28][3] , \memory[28][2] ,
         \memory[28][1] , \memory[28][0] , \memory[27][3] , \memory[27][2] ,
         \memory[27][1] , \memory[27][0] , \memory[26][3] , \memory[26][2] ,
         \memory[26][1] , \memory[26][0] , \memory[25][3] , \memory[25][2] ,
         \memory[25][1] , \memory[25][0] , \memory[24][3] , \memory[24][2] ,
         \memory[24][1] , \memory[24][0] , \memory[23][3] , \memory[23][2] ,
         \memory[23][1] , \memory[23][0] , \memory[22][3] , \memory[22][2] ,
         \memory[22][1] , \memory[22][0] , \memory[21][3] , \memory[21][2] ,
         \memory[21][1] , \memory[21][0] , \memory[20][3] , \memory[20][2] ,
         \memory[20][1] , \memory[20][0] , \memory[19][3] , \memory[19][2] ,
         \memory[19][1] , \memory[19][0] , \memory[18][3] , \memory[18][2] ,
         \memory[18][1] , \memory[18][0] , \memory[17][3] , \memory[17][2] ,
         \memory[17][1] , \memory[17][0] , \memory[16][3] , \memory[16][2] ,
         \memory[16][1] , \memory[16][0] , \memory[15][3] , \memory[15][2] ,
         \memory[15][1] , \memory[15][0] , \memory[14][3] , \memory[14][2] ,
         \memory[14][1] , \memory[14][0] , \memory[13][3] , \memory[13][2] ,
         \memory[13][1] , \memory[13][0] , \memory[12][3] , \memory[12][2] ,
         \memory[12][1] , \memory[12][0] , \memory[11][3] , \memory[11][2] ,
         \memory[11][1] , \memory[11][0] , \memory[10][3] , \memory[10][2] ,
         \memory[10][1] , \memory[10][0] , \memory[9][3] , \memory[9][2] ,
         \memory[9][1] , \memory[9][0] , \memory[8][3] , \memory[8][2] ,
         \memory[8][1] , \memory[8][0] , \memory[7][3] , \memory[7][2] ,
         \memory[7][1] , \memory[7][0] , \memory[6][3] , \memory[6][2] ,
         \memory[6][1] , \memory[6][0] , \memory[5][3] , \memory[5][2] ,
         \memory[5][1] , \memory[5][0] , \memory[4][3] , \memory[4][2] ,
         \memory[4][1] , \memory[4][0] , \memory[3][3] , \memory[3][2] ,
         \memory[3][1] , \memory[3][0] , \memory[2][3] , \memory[2][2] ,
         \memory[2][1] , \memory[2][0] , \memory[1][3] , \memory[1][2] ,
         \memory[1][1] , \memory[1][0] , \memory[0][3] , \memory[0][2] ,
         \memory[0][1] , \memory[0][0] , N61, N63, N65, N67, N69, N71, N73,
         N75, N77, N79, N81, N83, N85, N87, N89, N91, N93, N95, N97, N98, N99,
         N101, N103, N105, N107, N109, N111, N113, N115, N117, N119, N121,
         N123, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256,
         N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N282, N563, N564, N565, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582,
         N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593,
         N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604,
         N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615,
         N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648,
         N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659,
         N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670,
         N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681,
         N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692,
         N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703,
         N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714,
         N1035, N1037, N1039, N1041, N1043, N1045, N1047, N1049, N1051, N1053,
         N1055, N1057, N1059, N1061, N1063, N1065, N1067, N1069, N1071, N1073,
         N1075, N1077, N1079, N1081, N1083, N1085, N1087, N1089, N1091, N1093,
         N1095, N1097, N1099, N1101, N1103, N1105, N1107, N1109, N1111, N1113,
         N1115, N1117, N1119, N1121, N1123, N1125, N1127, N1129, N1131, N1133,
         N1135, N1137, N1139, N1141, N1143, N1145, N1147, N1149, N1151, N1153,
         N1155, N1157, N1159, N1161, N1163, N1165, N1167, N1169, N1171, N1173,
         N1175, N1177, N1179, N1181, N1183, N1185, N1187, N1189, N1191, N1193,
         N1195, N1197, N1199, N1201, N1203, N1205, N1207, N1209, N1211, N1213,
         N1215, N1217, N1219, N1221, N1223, N1225, N1227, N1229, N1231, N1233,
         N1235, N1237, N1239, N1241, N1243, N1245, N1247, N1249, N1251, N1253,
         N1255, N1257, N1259, N1261, N1263, N1265, N1267, N1269, N1271, N1273,
         N1275, N1277, N1279, N1281, N1283, N1285, N1291, N1293, N1295, N1297,
         N1299, N1301, N1303, N1305, N1307, N1309, N1311, N1313, N1315, N1317,
         N1319, N1321, N1323, N1325, N1327, N1329, N1331, N1333, N1335, N1337,
         N1339, N1341, N1343, N1345, N1347, N1349, N1351, N1482, N1483, N1519,
         N1523, N1527, N1531, N1535, N1539, N1543, N1547, N1551, N1555, N1559,
         N1563, N1567, N1571, N1575, N1579, N1583, N1587, N1591, N1595, N1599,
         N1603, N1607, N1611, N1615, N1619, N1623, N1627, N1631, N1635, N1639,
         N1643, N1647, N1651, N1654, N1656, N1667, N1669, N1672, N1674, N1678,
         N1680, N1682, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691,
         N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701,
         N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711,
         N1712, N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720, N1721,
         N1722, N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730, N1731,
         N1732, N1733, N1735, N1736, N1738, N1739, N1741, N1742, N1744, N1745,
         N1747, N1748, N1750, N1751, N1753, N1754, N1756, N1757, N1759, N1760,
         N1762, N1763, N1765, N1766, N1768, N1769, N1771, N1772, N1774, N1775,
         N1777, N1778, N1780, N1781, N1783, N1784, N1786, N1787, N1789, N1790,
         N1792, N1793, N1795, N1796, N1798, N1799, N1801, N1802, N1804, N1805,
         N1807, N1808, N1810, N1811, N1813, N1814, N1816, N1820, N1823, N1829,
         N1831, N1832, N1834, N1835, N1837, N1838, N1840, N1841, N1843, N1844,
         N1846, N1847, N1849, N1850, N1852, N1853, N1855, N1856, N1858, N1859,
         N1861, N1862, N1864, N1865, N1867, N1868, N1870, N1871, N1873, N1874,
         N1876, N1877, N1879, N1880, N1882, N1883, N1885, N1886, N1888, N1889,
         N1891, N1892, N1894, N1895, N1897, N1898, N1900, N1901, N1903, N1904,
         N1906, N1907, N1909, N1910, N1912, N1913, N1915, N1916, N1918, N1919,
         N1921, N1922, N1924, N1925, N1927, N1928, N1930, N1931, N1933, N1934,
         N1936, N1937, N1939, N1940, N1942, N1943, N1945, N1946, N1948, N1949,
         N1951, N1952, N1954, N1955, N1957, N1958, N1960, N1961, N1963, N1964,
         N1966, N1967, N1969, N1970, N1972, N1973, N1975, N1976, N1978, N1979,
         N1981, N1982, N1984, N1985, N1987, N1988, N1990, N1991, N1993, N1994,
         N1996, N1997, N1999, N2000, N2002, N2003, N2005, N2006, N2008, N2009,
         N2011, N2012, N2014, N2015, N2017, N2018, N2020, N2021, N2023, N2024,
         N2026, N2027, N2029, N2030, N2032, N2033, N2035, N2036, N2038, N2039,
         N2041, N2042, N2044, N2045, N2047, N2048, N2050, N2051, N2053, N2054,
         N2056, N2057, N2059, N2060, N2062, N2063, N2065, N2066, N2068, N2069,
         N2071, N2072, N2074, N2075, N2077, N2078, N2080, N2081, N2083, N2084,
         N2086, N2087, N2089, N2090, N2092, N2093, N2095, N2096, N2098, N2099,
         N2101, N2102, N2104, N2105, N2107, N2108, N2110, N2111, N2113, N2114,
         N2116, N2117, N2119, N2120, N2122, N2123, N2125, N2126, N2128, N2129,
         N2131, N2132, N2134, N2135, N2137, N2138, N2140, N2141, N2143, N2144,
         N2146, N2147, N2149, N2150, N2152, N2153, N2155, N2156, N2158, N2159,
         N2161, N2162, N2164, N2165, N2167, N2168, N2170, N2171, N2173, N2174,
         N2176, N2177, N2179, N2180, N2182, N2183, N2185, N2186, N2188, n12,
         n13, n14, n15, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690;
  wire   [31:0] counter;

  CAN2X2 C3473 ( .A(n672), .B(\memory[30][0] ), .Z(N2188) );
  CAN2X2 C3472 ( .A(n653), .B(\memory[31][0] ), .Z(N2186) );
  COR2X1 C3471 ( .A(N2186), .B(N2188), .Z(N714) );
  CAN2X2 C3469 ( .A(n663), .B(\memory[30][1] ), .Z(N2185) );
  CAN2X2 C3468 ( .A(n662), .B(\memory[31][1] ), .Z(N2183) );
  COR2X1 C3467 ( .A(N2183), .B(N2185), .Z(N713) );
  CAN2X2 C3465 ( .A(n672), .B(\memory[30][2] ), .Z(N2182) );
  CAN2X2 C3464 ( .A(n653), .B(\memory[31][2] ), .Z(N2180) );
  COR2X1 C3463 ( .A(N2180), .B(N2182), .Z(N712) );
  CAN2X2 C3461 ( .A(n663), .B(\memory[30][3] ), .Z(N2179) );
  CAN2X2 C3460 ( .A(n662), .B(\memory[31][3] ), .Z(N2177) );
  COR2X1 C3459 ( .A(N2177), .B(N2179), .Z(N711) );
  CAN2X2 C3457 ( .A(n671), .B(\memory[29][0] ), .Z(N2176) );
  CAN2X2 C3456 ( .A(n653), .B(\memory[30][0] ), .Z(N2174) );
  COR2X1 C3455 ( .A(N2174), .B(N2176), .Z(N710) );
  CAN2X2 C3453 ( .A(n663), .B(\memory[29][1] ), .Z(N2173) );
  CAN2X2 C3452 ( .A(n662), .B(\memory[30][1] ), .Z(N2171) );
  COR2X1 C3451 ( .A(N2171), .B(N2173), .Z(N709) );
  CAN2X2 C3449 ( .A(n672), .B(\memory[29][2] ), .Z(N2170) );
  CAN2X2 C3448 ( .A(n653), .B(\memory[30][2] ), .Z(N2168) );
  COR2X1 C3447 ( .A(N2168), .B(N2170), .Z(N708) );
  CAN2X2 C3445 ( .A(n663), .B(\memory[29][3] ), .Z(N2167) );
  CAN2X2 C3444 ( .A(n662), .B(\memory[30][3] ), .Z(N2165) );
  COR2X1 C3443 ( .A(N2165), .B(N2167), .Z(N707) );
  CAN2X2 C3441 ( .A(n671), .B(\memory[28][0] ), .Z(N2164) );
  CAN2X2 C3440 ( .A(n653), .B(\memory[29][0] ), .Z(N2162) );
  COR2X1 C3439 ( .A(N2162), .B(N2164), .Z(N706) );
  CAN2X2 C3437 ( .A(n663), .B(\memory[28][1] ), .Z(N2161) );
  CAN2X2 C3436 ( .A(n661), .B(\memory[29][1] ), .Z(N2159) );
  COR2X1 C3435 ( .A(N2159), .B(N2161), .Z(N705) );
  CAN2X2 C3433 ( .A(n671), .B(\memory[28][2] ), .Z(N2158) );
  CAN2X2 C3432 ( .A(n653), .B(\memory[29][2] ), .Z(N2156) );
  COR2X1 C3431 ( .A(N2156), .B(N2158), .Z(N704) );
  CAN2X2 C3429 ( .A(n663), .B(\memory[28][3] ), .Z(N2155) );
  CAN2X2 C3428 ( .A(n661), .B(\memory[29][3] ), .Z(N2153) );
  COR2X1 C3427 ( .A(N2153), .B(N2155), .Z(N703) );
  CAN2X2 C3425 ( .A(n671), .B(\memory[27][0] ), .Z(N2152) );
  CAN2X2 C3424 ( .A(n653), .B(\memory[28][0] ), .Z(N2150) );
  COR2X1 C3423 ( .A(N2150), .B(N2152), .Z(N702) );
  CAN2X2 C3421 ( .A(n663), .B(\memory[27][1] ), .Z(N2149) );
  CAN2X2 C3420 ( .A(n661), .B(\memory[28][1] ), .Z(N2147) );
  COR2X1 C3419 ( .A(N2147), .B(N2149), .Z(N701) );
  CAN2X2 C3417 ( .A(n671), .B(\memory[27][2] ), .Z(N2146) );
  CAN2X2 C3416 ( .A(n653), .B(\memory[28][2] ), .Z(N2144) );
  COR2X1 C3415 ( .A(N2144), .B(N2146), .Z(N700) );
  CAN2X2 C3413 ( .A(n663), .B(\memory[27][3] ), .Z(N2143) );
  CAN2X2 C3412 ( .A(n661), .B(\memory[28][3] ), .Z(N2141) );
  COR2X1 C3411 ( .A(N2141), .B(N2143), .Z(N699) );
  CAN2X2 C3409 ( .A(n671), .B(\memory[26][0] ), .Z(N2140) );
  CAN2X2 C3408 ( .A(n653), .B(\memory[27][0] ), .Z(N2138) );
  COR2X1 C3407 ( .A(N2138), .B(N2140), .Z(N698) );
  CAN2X2 C3405 ( .A(n663), .B(\memory[26][1] ), .Z(N2137) );
  CAN2X2 C3404 ( .A(n661), .B(\memory[27][1] ), .Z(N2135) );
  COR2X1 C3403 ( .A(N2135), .B(N2137), .Z(N697) );
  CAN2X2 C3401 ( .A(n671), .B(\memory[26][2] ), .Z(N2134) );
  CAN2X2 C3400 ( .A(n653), .B(\memory[27][2] ), .Z(N2132) );
  COR2X1 C3399 ( .A(N2132), .B(N2134), .Z(N696) );
  CAN2X2 C3397 ( .A(n663), .B(\memory[26][3] ), .Z(N2131) );
  CAN2X2 C3396 ( .A(n661), .B(\memory[27][3] ), .Z(N2129) );
  COR2X1 C3395 ( .A(N2129), .B(N2131), .Z(N695) );
  CAN2X2 C3393 ( .A(n671), .B(\memory[25][0] ), .Z(N2128) );
  CAN2X2 C3392 ( .A(n653), .B(\memory[26][0] ), .Z(N2126) );
  COR2X1 C3391 ( .A(N2126), .B(N2128), .Z(N694) );
  CAN2X2 C3389 ( .A(n663), .B(\memory[25][1] ), .Z(N2125) );
  CAN2X2 C3388 ( .A(n661), .B(\memory[26][1] ), .Z(N2123) );
  COR2X1 C3387 ( .A(N2123), .B(N2125), .Z(N693) );
  CAN2X2 C3385 ( .A(n671), .B(\memory[25][2] ), .Z(N2122) );
  CAN2X2 C3384 ( .A(n653), .B(\memory[26][2] ), .Z(N2120) );
  COR2X1 C3383 ( .A(N2120), .B(N2122), .Z(N692) );
  CAN2X2 C3381 ( .A(n663), .B(\memory[25][3] ), .Z(N2119) );
  CAN2X2 C3380 ( .A(n661), .B(\memory[26][3] ), .Z(N2117) );
  COR2X1 C3379 ( .A(N2117), .B(N2119), .Z(N691) );
  CAN2X2 C3377 ( .A(n671), .B(\memory[24][0] ), .Z(N2116) );
  CAN2X2 C3376 ( .A(n654), .B(\memory[25][0] ), .Z(N2114) );
  COR2X1 C3375 ( .A(N2114), .B(N2116), .Z(N690) );
  CAN2X2 C3373 ( .A(n664), .B(\memory[24][1] ), .Z(N2113) );
  CAN2X2 C3372 ( .A(n661), .B(\memory[25][1] ), .Z(N2111) );
  COR2X1 C3371 ( .A(N2111), .B(N2113), .Z(N689) );
  CAN2X2 C3369 ( .A(n671), .B(\memory[24][2] ), .Z(N2110) );
  CAN2X2 C3368 ( .A(n653), .B(\memory[25][2] ), .Z(N2108) );
  COR2X1 C3367 ( .A(N2108), .B(N2110), .Z(N688) );
  CAN2X2 C3365 ( .A(n663), .B(\memory[24][3] ), .Z(N2107) );
  CAN2X2 C3364 ( .A(n661), .B(\memory[25][3] ), .Z(N2105) );
  COR2X1 C3363 ( .A(N2105), .B(N2107), .Z(N687) );
  CAN2X2 C3361 ( .A(n671), .B(\memory[23][0] ), .Z(N2104) );
  CAN2X2 C3360 ( .A(n654), .B(\memory[24][0] ), .Z(N2102) );
  COR2X1 C3359 ( .A(N2102), .B(N2104), .Z(N686) );
  CAN2X2 C3357 ( .A(n664), .B(\memory[23][1] ), .Z(N2101) );
  CAN2X2 C3356 ( .A(n661), .B(\memory[24][1] ), .Z(N2099) );
  COR2X1 C3355 ( .A(N2099), .B(N2101), .Z(N685) );
  CAN2X2 C3353 ( .A(n671), .B(\memory[23][2] ), .Z(N2098) );
  CAN2X2 C3352 ( .A(n654), .B(\memory[24][2] ), .Z(N2096) );
  COR2X1 C3351 ( .A(N2096), .B(N2098), .Z(N684) );
  CAN2X2 C3349 ( .A(n664), .B(\memory[23][3] ), .Z(N2095) );
  CAN2X2 C3348 ( .A(n661), .B(\memory[24][3] ), .Z(N2093) );
  COR2X1 C3347 ( .A(N2093), .B(N2095), .Z(N683) );
  CAN2X2 C3345 ( .A(n670), .B(\memory[22][0] ), .Z(N2092) );
  CAN2X2 C3344 ( .A(n654), .B(\memory[23][0] ), .Z(N2090) );
  COR2X1 C3343 ( .A(N2090), .B(N2092), .Z(N682) );
  CAN2X2 C3341 ( .A(n664), .B(\memory[22][1] ), .Z(N2089) );
  CAN2X2 C3340 ( .A(n660), .B(\memory[23][1] ), .Z(N2087) );
  COR2X1 C3339 ( .A(N2087), .B(N2089), .Z(N681) );
  CAN2X2 C3337 ( .A(n670), .B(\memory[22][2] ), .Z(N2086) );
  CAN2X2 C3336 ( .A(n654), .B(\memory[23][2] ), .Z(N2084) );
  COR2X1 C3335 ( .A(N2084), .B(N2086), .Z(N680) );
  CAN2X2 C3333 ( .A(n664), .B(\memory[22][3] ), .Z(N2083) );
  CAN2X2 C3332 ( .A(n661), .B(\memory[23][3] ), .Z(N2081) );
  COR2X1 C3331 ( .A(N2081), .B(N2083), .Z(N679) );
  CAN2X2 C3329 ( .A(n670), .B(\memory[21][0] ), .Z(N2080) );
  CAN2X2 C3328 ( .A(n654), .B(\memory[22][0] ), .Z(N2078) );
  COR2X1 C3327 ( .A(N2078), .B(N2080), .Z(N678) );
  CAN2X2 C3325 ( .A(n664), .B(\memory[21][1] ), .Z(N2077) );
  CAN2X2 C3324 ( .A(n660), .B(\memory[22][1] ), .Z(N2075) );
  COR2X1 C3323 ( .A(N2075), .B(N2077), .Z(N677) );
  CAN2X2 C3321 ( .A(n670), .B(\memory[21][2] ), .Z(N2074) );
  CAN2X2 C3320 ( .A(n654), .B(\memory[22][2] ), .Z(N2072) );
  COR2X1 C3319 ( .A(N2072), .B(N2074), .Z(N676) );
  CAN2X2 C3317 ( .A(n664), .B(\memory[21][3] ), .Z(N2071) );
  CAN2X2 C3316 ( .A(n660), .B(\memory[22][3] ), .Z(N2069) );
  COR2X1 C3315 ( .A(N2069), .B(N2071), .Z(N675) );
  CAN2X2 C3313 ( .A(n670), .B(\memory[20][0] ), .Z(N2068) );
  CAN2X2 C3312 ( .A(n654), .B(\memory[21][0] ), .Z(N2066) );
  COR2X1 C3311 ( .A(N2066), .B(N2068), .Z(N674) );
  CAN2X2 C3309 ( .A(n664), .B(\memory[20][1] ), .Z(N2065) );
  CAN2X2 C3308 ( .A(n660), .B(\memory[21][1] ), .Z(N2063) );
  COR2X1 C3307 ( .A(N2063), .B(N2065), .Z(N673) );
  CAN2X2 C3305 ( .A(n670), .B(\memory[20][2] ), .Z(N2062) );
  CAN2X2 C3304 ( .A(n654), .B(\memory[21][2] ), .Z(N2060) );
  COR2X1 C3303 ( .A(N2060), .B(N2062), .Z(N672) );
  CAN2X2 C3301 ( .A(n664), .B(\memory[20][3] ), .Z(N2059) );
  CAN2X2 C3300 ( .A(n660), .B(\memory[21][3] ), .Z(N2057) );
  COR2X1 C3299 ( .A(N2057), .B(N2059), .Z(N671) );
  CAN2X2 C3297 ( .A(n670), .B(\memory[19][0] ), .Z(N2056) );
  CAN2X2 C3296 ( .A(n654), .B(\memory[20][0] ), .Z(N2054) );
  COR2X1 C3295 ( .A(N2054), .B(N2056), .Z(N670) );
  CAN2X2 C3293 ( .A(n664), .B(\memory[19][1] ), .Z(N2053) );
  CAN2X2 C3292 ( .A(n660), .B(\memory[20][1] ), .Z(N2051) );
  COR2X1 C3291 ( .A(N2051), .B(N2053), .Z(N669) );
  CAN2X2 C3289 ( .A(n670), .B(\memory[19][2] ), .Z(N2050) );
  CAN2X2 C3288 ( .A(n654), .B(\memory[20][2] ), .Z(N2048) );
  COR2X1 C3287 ( .A(N2048), .B(N2050), .Z(N668) );
  CAN2X2 C3285 ( .A(n664), .B(\memory[19][3] ), .Z(N2047) );
  CAN2X2 C3284 ( .A(n660), .B(\memory[20][3] ), .Z(N2045) );
  COR2X1 C3283 ( .A(N2045), .B(N2047), .Z(N667) );
  CAN2X2 C3281 ( .A(n670), .B(\memory[18][0] ), .Z(N2044) );
  CAN2X2 C3280 ( .A(n654), .B(\memory[19][0] ), .Z(N2042) );
  COR2X1 C3279 ( .A(N2042), .B(N2044), .Z(N666) );
  CAN2X2 C3277 ( .A(n664), .B(\memory[18][1] ), .Z(N2041) );
  CAN2X2 C3276 ( .A(n660), .B(\memory[19][1] ), .Z(N2039) );
  COR2X1 C3275 ( .A(N2039), .B(N2041), .Z(N665) );
  CAN2X2 C3273 ( .A(n670), .B(\memory[18][2] ), .Z(N2038) );
  CAN2X2 C3272 ( .A(n654), .B(\memory[19][2] ), .Z(N2036) );
  COR2X1 C3271 ( .A(N2036), .B(N2038), .Z(N664) );
  CAN2X2 C3269 ( .A(n664), .B(\memory[18][3] ), .Z(N2035) );
  CAN2X2 C3268 ( .A(n660), .B(\memory[19][3] ), .Z(N2033) );
  COR2X1 C3267 ( .A(N2033), .B(N2035), .Z(N663) );
  CAN2X2 C3265 ( .A(n670), .B(\memory[17][0] ), .Z(N2032) );
  CAN2X2 C3264 ( .A(n655), .B(\memory[18][0] ), .Z(N2030) );
  COR2X1 C3263 ( .A(N2030), .B(N2032), .Z(N662) );
  CAN2X2 C3261 ( .A(n665), .B(\memory[17][1] ), .Z(N2029) );
  CAN2X2 C3260 ( .A(n660), .B(\memory[18][1] ), .Z(N2027) );
  COR2X1 C3259 ( .A(N2027), .B(N2029), .Z(N661) );
  CAN2X2 C3257 ( .A(n670), .B(\memory[17][2] ), .Z(N2026) );
  CAN2X2 C3256 ( .A(n655), .B(\memory[18][2] ), .Z(N2024) );
  COR2X1 C3255 ( .A(N2024), .B(N2026), .Z(N660) );
  CAN2X2 C3253 ( .A(n665), .B(\memory[17][3] ), .Z(N2023) );
  CAN2X2 C3252 ( .A(n660), .B(\memory[18][3] ), .Z(N2021) );
  COR2X1 C3251 ( .A(N2021), .B(N2023), .Z(N659) );
  CAN2X2 C3249 ( .A(n669), .B(\memory[16][0] ), .Z(N2020) );
  CAN2X2 C3248 ( .A(n655), .B(\memory[17][0] ), .Z(N2018) );
  COR2X1 C3247 ( .A(N2018), .B(N2020), .Z(N658) );
  CAN2X2 C3245 ( .A(n665), .B(\memory[16][1] ), .Z(N2017) );
  CAN2X2 C3244 ( .A(n660), .B(\memory[17][1] ), .Z(N2015) );
  COR2X1 C3243 ( .A(N2015), .B(N2017), .Z(N657) );
  CAN2X2 C3241 ( .A(n670), .B(\memory[16][2] ), .Z(N2014) );
  CAN2X2 C3240 ( .A(n655), .B(\memory[17][2] ), .Z(N2012) );
  COR2X1 C3239 ( .A(N2012), .B(N2014), .Z(N656) );
  CAN2X2 C3237 ( .A(n665), .B(\memory[16][3] ), .Z(N2011) );
  CAN2X2 C3236 ( .A(n660), .B(\memory[17][3] ), .Z(N2009) );
  COR2X1 C3235 ( .A(N2009), .B(N2011), .Z(N655) );
  CAN2X2 C3233 ( .A(n669), .B(\memory[15][0] ), .Z(N2008) );
  CAN2X2 C3232 ( .A(n655), .B(\memory[16][0] ), .Z(N2006) );
  COR2X1 C3231 ( .A(N2006), .B(N2008), .Z(N654) );
  CAN2X2 C3229 ( .A(n665), .B(\memory[15][1] ), .Z(N2005) );
  CAN2X2 C3228 ( .A(n659), .B(\memory[16][1] ), .Z(N2003) );
  COR2X1 C3227 ( .A(N2003), .B(N2005), .Z(N653) );
  CAN2X2 C3225 ( .A(n669), .B(\memory[15][2] ), .Z(N2002) );
  CAN2X2 C3224 ( .A(n655), .B(\memory[16][2] ), .Z(N2000) );
  COR2X1 C3223 ( .A(N2000), .B(N2002), .Z(N652) );
  CAN2X2 C3221 ( .A(n665), .B(\memory[15][3] ), .Z(N1999) );
  CAN2X2 C3220 ( .A(n659), .B(\memory[16][3] ), .Z(N1997) );
  COR2X1 C3219 ( .A(N1997), .B(N1999), .Z(N651) );
  CAN2X2 C3217 ( .A(n669), .B(\memory[14][0] ), .Z(N1996) );
  CAN2X2 C3216 ( .A(n655), .B(\memory[15][0] ), .Z(N1994) );
  COR2X1 C3215 ( .A(N1994), .B(N1996), .Z(N650) );
  CAN2X2 C3213 ( .A(n665), .B(\memory[14][1] ), .Z(N1993) );
  CAN2X2 C3212 ( .A(n659), .B(\memory[15][1] ), .Z(N1991) );
  COR2X1 C3211 ( .A(N1991), .B(N1993), .Z(N649) );
  CAN2X2 C3209 ( .A(n669), .B(\memory[14][2] ), .Z(N1990) );
  CAN2X2 C3208 ( .A(n655), .B(\memory[15][2] ), .Z(N1988) );
  COR2X1 C3207 ( .A(N1988), .B(N1990), .Z(N648) );
  CAN2X2 C3205 ( .A(n665), .B(\memory[14][3] ), .Z(N1987) );
  CAN2X2 C3204 ( .A(n659), .B(\memory[15][3] ), .Z(N1985) );
  COR2X1 C3203 ( .A(N1985), .B(N1987), .Z(N647) );
  CAN2X2 C3201 ( .A(n669), .B(\memory[13][0] ), .Z(N1984) );
  CAN2X2 C3200 ( .A(n655), .B(\memory[14][0] ), .Z(N1982) );
  COR2X1 C3199 ( .A(N1982), .B(N1984), .Z(N646) );
  CAN2X2 C3197 ( .A(n665), .B(\memory[13][1] ), .Z(N1981) );
  CAN2X2 C3196 ( .A(n659), .B(\memory[14][1] ), .Z(N1979) );
  COR2X1 C3195 ( .A(N1979), .B(N1981), .Z(N645) );
  CAN2X2 C3193 ( .A(n669), .B(\memory[13][2] ), .Z(N1978) );
  CAN2X2 C3192 ( .A(n655), .B(\memory[14][2] ), .Z(N1976) );
  COR2X1 C3191 ( .A(N1976), .B(N1978), .Z(N644) );
  CAN2X2 C3189 ( .A(n665), .B(\memory[13][3] ), .Z(N1975) );
  CAN2X2 C3188 ( .A(n659), .B(\memory[14][3] ), .Z(N1973) );
  COR2X1 C3187 ( .A(N1973), .B(N1975), .Z(N643) );
  CAN2X2 C3185 ( .A(n669), .B(\memory[12][0] ), .Z(N1972) );
  CAN2X2 C3184 ( .A(n655), .B(\memory[13][0] ), .Z(N1970) );
  COR2X1 C3183 ( .A(N1970), .B(N1972), .Z(N642) );
  CAN2X2 C3181 ( .A(n665), .B(\memory[12][1] ), .Z(N1969) );
  CAN2X2 C3180 ( .A(n659), .B(\memory[13][1] ), .Z(N1967) );
  COR2X1 C3179 ( .A(N1967), .B(N1969), .Z(N641) );
  CAN2X2 C3177 ( .A(n669), .B(\memory[12][2] ), .Z(N1966) );
  CAN2X2 C3176 ( .A(n655), .B(\memory[13][2] ), .Z(N1964) );
  COR2X1 C3175 ( .A(N1964), .B(N1966), .Z(N640) );
  CAN2X2 C3173 ( .A(n665), .B(\memory[12][3] ), .Z(N1963) );
  CAN2X2 C3172 ( .A(n659), .B(\memory[13][3] ), .Z(N1961) );
  COR2X1 C3171 ( .A(N1961), .B(N1963), .Z(N639) );
  CAN2X2 C3169 ( .A(n669), .B(\memory[11][0] ), .Z(N1960) );
  CAN2X2 C3168 ( .A(n656), .B(\memory[12][0] ), .Z(N1958) );
  COR2X1 C3167 ( .A(N1958), .B(N1960), .Z(N638) );
  CAN2X2 C3165 ( .A(n666), .B(\memory[11][1] ), .Z(N1957) );
  CAN2X2 C3164 ( .A(n659), .B(\memory[12][1] ), .Z(N1955) );
  COR2X1 C3163 ( .A(N1955), .B(N1957), .Z(N637) );
  CAN2X2 C3161 ( .A(n669), .B(\memory[11][2] ), .Z(N1954) );
  CAN2X2 C3160 ( .A(n655), .B(\memory[12][2] ), .Z(N1952) );
  COR2X1 C3159 ( .A(N1952), .B(N1954), .Z(N636) );
  CAN2X2 C3157 ( .A(n665), .B(\memory[11][3] ), .Z(N1951) );
  CAN2X2 C3156 ( .A(n659), .B(\memory[12][3] ), .Z(N1949) );
  COR2X1 C3155 ( .A(N1949), .B(N1951), .Z(N635) );
  CAN2X2 C3153 ( .A(n669), .B(\memory[10][0] ), .Z(N1948) );
  CAN2X2 C3152 ( .A(n656), .B(\memory[11][0] ), .Z(N1946) );
  COR2X1 C3151 ( .A(N1946), .B(N1948), .Z(N634) );
  CAN2X2 C3149 ( .A(n666), .B(\memory[10][1] ), .Z(N1945) );
  CAN2X2 C3148 ( .A(n659), .B(\memory[11][1] ), .Z(N1943) );
  COR2X1 C3147 ( .A(N1943), .B(N1945), .Z(N633) );
  CAN2X2 C3145 ( .A(n669), .B(\memory[10][2] ), .Z(N1942) );
  CAN2X2 C3144 ( .A(n656), .B(\memory[11][2] ), .Z(N1940) );
  COR2X1 C3143 ( .A(N1940), .B(N1942), .Z(N632) );
  CAN2X2 C3141 ( .A(n666), .B(\memory[10][3] ), .Z(N1939) );
  CAN2X2 C3140 ( .A(n659), .B(\memory[11][3] ), .Z(N1937) );
  COR2X1 C3139 ( .A(N1937), .B(N1939), .Z(N631) );
  CAN2X2 C3137 ( .A(n668), .B(\memory[9][0] ), .Z(N1936) );
  CAN2X2 C3136 ( .A(n656), .B(\memory[10][0] ), .Z(N1934) );
  COR2X1 C3135 ( .A(N1934), .B(N1936), .Z(N630) );
  CAN2X2 C3133 ( .A(n666), .B(\memory[9][1] ), .Z(N1933) );
  CAN2X2 C3132 ( .A(n658), .B(\memory[10][1] ), .Z(N1931) );
  COR2X1 C3131 ( .A(N1931), .B(N1933), .Z(N629) );
  CAN2X2 C3129 ( .A(n668), .B(\memory[9][2] ), .Z(N1930) );
  CAN2X2 C3128 ( .A(n656), .B(\memory[10][2] ), .Z(N1928) );
  COR2X1 C3127 ( .A(N1928), .B(N1930), .Z(N628) );
  CAN2X2 C3125 ( .A(n666), .B(\memory[9][3] ), .Z(N1927) );
  CAN2X2 C3124 ( .A(n659), .B(\memory[10][3] ), .Z(N1925) );
  COR2X1 C3123 ( .A(N1925), .B(N1927), .Z(N627) );
  CAN2X2 C3121 ( .A(n668), .B(\memory[8][0] ), .Z(N1924) );
  CAN2X2 C3120 ( .A(n656), .B(\memory[9][0] ), .Z(N1922) );
  COR2X1 C3119 ( .A(N1922), .B(N1924), .Z(N626) );
  CAN2X2 C3117 ( .A(n666), .B(\memory[8][1] ), .Z(N1921) );
  CAN2X2 C3116 ( .A(n658), .B(\memory[9][1] ), .Z(N1919) );
  COR2X1 C3115 ( .A(N1919), .B(N1921), .Z(N625) );
  CAN2X2 C3113 ( .A(n668), .B(\memory[8][2] ), .Z(N1918) );
  CAN2X2 C3112 ( .A(n656), .B(\memory[9][2] ), .Z(N1916) );
  COR2X1 C3111 ( .A(N1916), .B(N1918), .Z(N624) );
  CAN2X2 C3109 ( .A(n666), .B(\memory[8][3] ), .Z(N1915) );
  CAN2X2 C3108 ( .A(n658), .B(\memory[9][3] ), .Z(N1913) );
  COR2X1 C3107 ( .A(N1913), .B(N1915), .Z(N623) );
  CAN2X2 C3105 ( .A(n668), .B(\memory[7][0] ), .Z(N1912) );
  CAN2X2 C3104 ( .A(n656), .B(\memory[8][0] ), .Z(N1910) );
  COR2X1 C3103 ( .A(N1910), .B(N1912), .Z(N622) );
  CAN2X2 C3101 ( .A(n666), .B(\memory[7][1] ), .Z(N1909) );
  CAN2X2 C3100 ( .A(n658), .B(\memory[8][1] ), .Z(N1907) );
  COR2X1 C3099 ( .A(N1907), .B(N1909), .Z(N621) );
  CAN2X2 C3097 ( .A(n668), .B(\memory[7][2] ), .Z(N1906) );
  CAN2X2 C3096 ( .A(n656), .B(\memory[8][2] ), .Z(N1904) );
  COR2X1 C3095 ( .A(N1904), .B(N1906), .Z(N620) );
  CAN2X2 C3093 ( .A(n666), .B(\memory[7][3] ), .Z(N1903) );
  CAN2X2 C3092 ( .A(n658), .B(\memory[8][3] ), .Z(N1901) );
  COR2X1 C3091 ( .A(N1901), .B(N1903), .Z(N619) );
  CAN2X2 C3089 ( .A(n668), .B(\memory[6][0] ), .Z(N1900) );
  CAN2X2 C3088 ( .A(n656), .B(\memory[7][0] ), .Z(N1898) );
  COR2X1 C3087 ( .A(N1898), .B(N1900), .Z(N618) );
  CAN2X2 C3085 ( .A(n666), .B(\memory[6][1] ), .Z(N1897) );
  CAN2X2 C3084 ( .A(n658), .B(\memory[7][1] ), .Z(N1895) );
  COR2X1 C3083 ( .A(N1895), .B(N1897), .Z(N617) );
  CAN2X2 C3081 ( .A(n668), .B(\memory[6][2] ), .Z(N1894) );
  CAN2X2 C3080 ( .A(n656), .B(\memory[7][2] ), .Z(N1892) );
  COR2X1 C3079 ( .A(N1892), .B(N1894), .Z(N616) );
  CAN2X2 C3077 ( .A(n666), .B(\memory[6][3] ), .Z(N1891) );
  CAN2X2 C3076 ( .A(n658), .B(\memory[7][3] ), .Z(N1889) );
  COR2X1 C3075 ( .A(N1889), .B(N1891), .Z(N615) );
  CAN2X2 C3073 ( .A(n668), .B(\memory[5][0] ), .Z(N1888) );
  CAN2X2 C3072 ( .A(n656), .B(\memory[6][0] ), .Z(N1886) );
  COR2X1 C3071 ( .A(N1886), .B(N1888), .Z(N614) );
  CAN2X2 C3069 ( .A(n666), .B(\memory[5][1] ), .Z(N1885) );
  CAN2X2 C3068 ( .A(n658), .B(\memory[6][1] ), .Z(N1883) );
  COR2X1 C3067 ( .A(N1883), .B(N1885), .Z(N613) );
  CAN2X2 C3065 ( .A(n668), .B(\memory[5][2] ), .Z(N1882) );
  CAN2X2 C3064 ( .A(n656), .B(\memory[6][2] ), .Z(N1880) );
  COR2X1 C3063 ( .A(N1880), .B(N1882), .Z(N612) );
  CAN2X2 C3061 ( .A(n666), .B(\memory[5][3] ), .Z(N1879) );
  CAN2X2 C3060 ( .A(n658), .B(\memory[6][3] ), .Z(N1877) );
  COR2X1 C3059 ( .A(N1877), .B(N1879), .Z(N611) );
  CAN2X2 C3057 ( .A(n668), .B(\memory[4][0] ), .Z(N1876) );
  CAN2X2 C3056 ( .A(n657), .B(\memory[5][0] ), .Z(N1874) );
  COR2X1 C3055 ( .A(N1874), .B(N1876), .Z(N610) );
  CAN2X2 C3053 ( .A(n667), .B(\memory[4][1] ), .Z(N1873) );
  CAN2X2 C3052 ( .A(n658), .B(\memory[5][1] ), .Z(N1871) );
  COR2X1 C3051 ( .A(N1871), .B(N1873), .Z(N609) );
  CAN2X2 C3049 ( .A(n668), .B(\memory[4][2] ), .Z(N1870) );
  CAN2X2 C3048 ( .A(n657), .B(\memory[5][2] ), .Z(N1868) );
  COR2X1 C3047 ( .A(N1868), .B(N1870), .Z(N608) );
  CAN2X2 C3045 ( .A(n667), .B(\memory[4][3] ), .Z(N1867) );
  CAN2X2 C3044 ( .A(n658), .B(\memory[5][3] ), .Z(N1865) );
  COR2X1 C3043 ( .A(N1865), .B(N1867), .Z(N607) );
  CAN2X2 C3041 ( .A(n667), .B(\memory[3][0] ), .Z(N1864) );
  CAN2X2 C3040 ( .A(n657), .B(\memory[4][0] ), .Z(N1862) );
  COR2X1 C3039 ( .A(N1862), .B(N1864), .Z(N606) );
  CAN2X2 C3037 ( .A(n667), .B(\memory[3][1] ), .Z(N1861) );
  CAN2X2 C3036 ( .A(n658), .B(\memory[4][1] ), .Z(N1859) );
  COR2X1 C3035 ( .A(N1859), .B(N1861), .Z(N605) );
  CAN2X2 C3033 ( .A(n668), .B(\memory[3][2] ), .Z(N1858) );
  CAN2X2 C3032 ( .A(n657), .B(\memory[4][2] ), .Z(N1856) );
  COR2X1 C3031 ( .A(N1856), .B(N1858), .Z(N604) );
  CAN2X2 C3029 ( .A(n667), .B(\memory[3][3] ), .Z(N1855) );
  CAN2X2 C3028 ( .A(n658), .B(\memory[4][3] ), .Z(N1853) );
  COR2X1 C3027 ( .A(N1853), .B(N1855), .Z(N603) );
  CAN2X2 C3025 ( .A(n667), .B(\memory[2][0] ), .Z(N1852) );
  CAN2X2 C3024 ( .A(n657), .B(\memory[3][0] ), .Z(N1850) );
  COR2X1 C3023 ( .A(N1850), .B(N1852), .Z(N602) );
  CAN2X2 C3021 ( .A(n667), .B(\memory[2][1] ), .Z(N1849) );
  CAN2X2 C3020 ( .A(n657), .B(\memory[3][1] ), .Z(N1847) );
  COR2X1 C3019 ( .A(N1847), .B(N1849), .Z(N601) );
  CAN2X2 C3017 ( .A(n667), .B(\memory[2][2] ), .Z(N1846) );
  CAN2X2 C3016 ( .A(n657), .B(\memory[3][2] ), .Z(N1844) );
  COR2X1 C3015 ( .A(N1844), .B(N1846), .Z(N600) );
  CAN2X2 C3013 ( .A(n667), .B(\memory[2][3] ), .Z(N1843) );
  CAN2X2 C3012 ( .A(n657), .B(\memory[3][3] ), .Z(N1841) );
  COR2X1 C3011 ( .A(N1841), .B(N1843), .Z(N599) );
  CAN2X2 C3009 ( .A(n667), .B(\memory[1][0] ), .Z(N1840) );
  CAN2X2 C3008 ( .A(n657), .B(\memory[2][0] ), .Z(N1838) );
  COR2X1 C3007 ( .A(N1838), .B(N1840), .Z(N598) );
  CAN2X2 C3005 ( .A(n667), .B(\memory[1][1] ), .Z(N1837) );
  CAN2X2 C3004 ( .A(n657), .B(\memory[2][1] ), .Z(N1835) );
  COR2X1 C3003 ( .A(N1835), .B(N1837), .Z(N597) );
  CAN2X2 C3001 ( .A(n667), .B(\memory[1][2] ), .Z(N1834) );
  CAN2X2 C3000 ( .A(n657), .B(\memory[2][2] ), .Z(N1832) );
  COR2X1 C2999 ( .A(N1832), .B(N1834), .Z(N596) );
  CAN2X2 C2997 ( .A(n667), .B(\memory[1][3] ), .Z(N1831) );
  CAN2X2 C2996 ( .A(n657), .B(\memory[2][3] ), .Z(N1829) );
  COR2X1 C2995 ( .A(N1829), .B(N1831), .Z(N595) );
  CAN2X2 C2918 ( .A(n565), .B(N63), .Z(N1823) );
  CAN2X2 C2914 ( .A(n566), .B(N65), .Z(N1820) );
  CAN2X2 C2907 ( .A(n576), .B(counter[4]), .Z(N1816) );
  CAN2X2 C2906 ( .A(n568), .B(N69), .Z(N1814) );
  COR2X1 C2905 ( .A(N1814), .B(N1816), .Z(N275) );
  CAN2X2 C2903 ( .A(n577), .B(counter[5]), .Z(N1813) );
  CAN2X2 C2902 ( .A(n569), .B(N71), .Z(N1811) );
  COR2X1 C2901 ( .A(N1811), .B(N1813), .Z(N274) );
  CAN2X2 C2898 ( .A(n570), .B(N73), .Z(N1808) );
  COR2X1 C2897 ( .A(N1808), .B(N1810), .Z(N273) );
  CAN2X2 C2895 ( .A(n579), .B(counter[7]), .Z(N1807) );
  CAN2X2 C2894 ( .A(n571), .B(N75), .Z(N1805) );
  COR2X1 C2893 ( .A(N1805), .B(N1807), .Z(N272) );
  CAN2X2 C2891 ( .A(n596), .B(counter[8]), .Z(N1804) );
  CAN2X2 C2890 ( .A(n587), .B(N77), .Z(N1802) );
  COR2X1 C2889 ( .A(N1802), .B(N1804), .Z(N271) );
  CAN2X2 C2887 ( .A(n580), .B(counter[9]), .Z(N1801) );
  CAN2X2 C2886 ( .A(n572), .B(N79), .Z(N1799) );
  COR2X1 C2885 ( .A(N1799), .B(N1801), .Z(N270) );
  CAN2X2 C2883 ( .A(n597), .B(counter[10]), .Z(N1798) );
  CAN2X2 C2882 ( .A(n588), .B(N81), .Z(N1796) );
  COR2X1 C2881 ( .A(N1796), .B(N1798), .Z(N269) );
  CAN2X2 C2879 ( .A(n598), .B(counter[11]), .Z(N1795) );
  CAN2X2 C2878 ( .A(n589), .B(N83), .Z(N1793) );
  COR2X1 C2877 ( .A(N1793), .B(N1795), .Z(N268) );
  CAN2X2 C2875 ( .A(n599), .B(counter[12]), .Z(N1792) );
  CAN2X2 C2874 ( .A(n590), .B(N85), .Z(N1790) );
  COR2X1 C2873 ( .A(N1790), .B(N1792), .Z(N267) );
  CAN2X2 C2871 ( .A(n600), .B(counter[13]), .Z(N1789) );
  CAN2X2 C2870 ( .A(n591), .B(N87), .Z(N1787) );
  COR2X1 C2869 ( .A(N1787), .B(N1789), .Z(N266) );
  CAN2X2 C2867 ( .A(n601), .B(counter[14]), .Z(N1786) );
  CAN2X2 C2866 ( .A(n592), .B(N89), .Z(N1784) );
  COR2X1 C2865 ( .A(N1784), .B(N1786), .Z(N265) );
  CAN2X2 C2863 ( .A(n602), .B(counter[15]), .Z(N1783) );
  CAN2X2 C2862 ( .A(n593), .B(N91), .Z(N1781) );
  COR2X1 C2861 ( .A(N1781), .B(N1783), .Z(N264) );
  CAN2X2 C2859 ( .A(n603), .B(counter[16]), .Z(N1780) );
  CAN2X2 C2858 ( .A(n594), .B(N93), .Z(N1778) );
  COR2X1 C2857 ( .A(N1778), .B(N1780), .Z(N263) );
  CAN2X2 C2855 ( .A(n604), .B(counter[17]), .Z(N1777) );
  CAN2X2 C2854 ( .A(n595), .B(N95), .Z(N1775) );
  COR2X1 C2853 ( .A(N1775), .B(N1777), .Z(N262) );
  CAN2X2 C2850 ( .A(n565), .B(N97), .Z(N1772) );
  COR2X1 C2849 ( .A(N1772), .B(N1774), .Z(N261) );
  CAN2X2 C2847 ( .A(n580), .B(counter[19]), .Z(N1771) );
  CAN2X2 C2846 ( .A(n569), .B(N99), .Z(N1769) );
  COR2X1 C2845 ( .A(N1769), .B(N1771), .Z(N260) );
  CAN2X2 C2843 ( .A(n604), .B(counter[20]), .Z(N1768) );
  CAN2X2 C2842 ( .A(n564), .B(N101), .Z(N1766) );
  COR2X1 C2841 ( .A(N1766), .B(N1768), .Z(N259) );
  CAN2X2 C2838 ( .A(n567), .B(N103), .Z(N1763) );
  COR2X1 C2837 ( .A(N1763), .B(N1765), .Z(N258) );
  CAN2X2 C2834 ( .A(n566), .B(N105), .Z(N1760) );
  COR2X1 C2833 ( .A(N1760), .B(N1762), .Z(N257) );
  CAN2X2 C2830 ( .A(n590), .B(N107), .Z(N1757) );
  COR2X1 C2829 ( .A(N1757), .B(N1759), .Z(N256) );
  CAN2X2 C2826 ( .A(n588), .B(N109), .Z(N1754) );
  COR2X1 C2825 ( .A(N1754), .B(N1756), .Z(N255) );
  CAN2X2 C2822 ( .A(n587), .B(N111), .Z(N1751) );
  COR2X1 C2821 ( .A(N1751), .B(N1753), .Z(N254) );
  COR2X1 C2817 ( .A(N1748), .B(N1750), .Z(N253) );
  CAN2X2 C2815 ( .A(n578), .B(counter[27]), .Z(N1747) );
  COR2X1 C2813 ( .A(N1745), .B(N1747), .Z(N252) );
  CAN2X2 C2811 ( .A(n596), .B(counter[28]), .Z(N1744) );
  COR2X1 C2809 ( .A(N1742), .B(N1744), .Z(N251) );
  CAN2X2 C2806 ( .A(n570), .B(N119), .Z(N1739) );
  COR2X1 C2805 ( .A(N1739), .B(N1741), .Z(N250) );
  COR2X1 C2801 ( .A(N1736), .B(N1738), .Z(N249) );
  CAN2X2 C2798 ( .A(n591), .B(N123), .Z(N1733) );
  COR2X1 C2797 ( .A(N1733), .B(N1735), .Z(N248) );
  CAN2X2 C2689 ( .A(N1687), .B(N1700), .Z(N1732) );
  CAN2X2 C2688 ( .A(N1687), .B(N1699), .Z(N1731) );
  CAN2X2 C2687 ( .A(N1687), .B(N1698), .Z(N1730) );
  CAN2X2 C2686 ( .A(N1687), .B(N1697), .Z(N1729) );
  CAN2X2 C2685 ( .A(N1687), .B(N1696), .Z(N1728) );
  CAN2X2 C2684 ( .A(N1687), .B(N1695), .Z(N1727) );
  CAN2X2 C2683 ( .A(N1687), .B(N1694), .Z(N1726) );
  CAN2X2 C2682 ( .A(N1687), .B(N1693), .Z(N1725) );
  CAN2X2 C2681 ( .A(N1686), .B(N1700), .Z(N1724) );
  CAN2X2 C2680 ( .A(N1686), .B(N1699), .Z(N1723) );
  CAN2X2 C2679 ( .A(N1686), .B(N1698), .Z(N1722) );
  CAN2X2 C2678 ( .A(N1686), .B(N1697), .Z(N1721) );
  CAN2X2 C2677 ( .A(N1686), .B(N1696), .Z(N1720) );
  CAN2X2 C2676 ( .A(N1686), .B(N1695), .Z(N1719) );
  CAN2X2 C2675 ( .A(N1686), .B(N1694), .Z(N1718) );
  CAN2X2 C2674 ( .A(N1686), .B(N1693), .Z(N1717) );
  CAN2X2 C2673 ( .A(N1685), .B(N1700), .Z(N1716) );
  CAN2X2 C2672 ( .A(N1685), .B(N1699), .Z(N1715) );
  CAN2X2 C2671 ( .A(N1685), .B(N1698), .Z(N1714) );
  CAN2X2 C2670 ( .A(N1685), .B(N1697), .Z(N1713) );
  CAN2X2 C2669 ( .A(N1685), .B(N1696), .Z(N1712) );
  CAN2X2 C2668 ( .A(N1685), .B(N1695), .Z(N1711) );
  CAN2X2 C2667 ( .A(N1685), .B(N1694), .Z(N1710) );
  CAN2X2 C2666 ( .A(N1685), .B(N1693), .Z(N1709) );
  CAN2X2 C2665 ( .A(N1684), .B(N1700), .Z(N1708) );
  CAN2X2 C2664 ( .A(N1684), .B(N1699), .Z(N1707) );
  CAN2X2 C2663 ( .A(N1684), .B(N1698), .Z(N1706) );
  CAN2X2 C2662 ( .A(N1684), .B(N1697), .Z(N1705) );
  CAN2X2 C2661 ( .A(N1684), .B(N1696), .Z(N1704) );
  CAN2X2 C2660 ( .A(N1684), .B(N1695), .Z(N1703) );
  CAN2X2 C2659 ( .A(N1684), .B(N1694), .Z(N1702) );
  CAN2X2 C2658 ( .A(N1684), .B(N1693), .Z(N1701) );
  CAN2X2 C2657 ( .A(N1688), .B(N1692), .Z(N1700) );
  CAN2X2 C2656 ( .A(N1688), .B(N1691), .Z(N1699) );
  CAN2X2 C2655 ( .A(N1688), .B(N1690), .Z(N1698) );
  CAN2X2 C2654 ( .A(N1688), .B(N1689), .Z(N1697) );
  CIVX2 I_4 ( .A(N275), .Z(N3) );
  CIVX2 I_2 ( .A(N275), .Z(N1) );
  CFD1QX1 \memory_reg[30][3]  ( .D(n354), .CP(clock), .Q(\memory[30][3] ) );
  CFD1QX1 \memory_reg[30][1]  ( .D(n356), .CP(clock), .Q(\memory[30][1] ) );
  CFD1QX1 \memory_reg[0][1]  ( .D(n479), .CP(clock), .Q(\memory[0][1] ) );
  CFD4QXL empty_reg ( .D(n353), .CP(clock), .SD(reset), .Q(empty) );
  CAOR2X1 U3 ( .A(n652), .B(reset), .C(N1701), .D(n12), .Z(N1647) );
  CAOR1X1 U4 ( .A(n12), .B(N1702), .C(N1483), .Z(N1643) );
  CAOR1X1 U10 ( .A(n12), .B(N1703), .C(N1483), .Z(N1639) );
  CAOR1X1 U11 ( .A(n12), .B(N1704), .C(N1483), .Z(N1635) );
  CAOR1X1 U12 ( .A(n12), .B(N1705), .C(N1483), .Z(N1631) );
  CAOR1X1 U13 ( .A(n12), .B(N1706), .C(N1483), .Z(N1627) );
  CAOR1X1 U14 ( .A(n12), .B(N1707), .C(N1483), .Z(N1623) );
  CAOR1X1 U15 ( .A(n12), .B(N1708), .C(N1483), .Z(N1619) );
  CAOR1X1 U16 ( .A(n12), .B(N1709), .C(N1483), .Z(N1615) );
  CAOR1X1 U17 ( .A(n12), .B(N1710), .C(N1483), .Z(N1611) );
  CAOR1X1 U18 ( .A(n12), .B(N1711), .C(N1483), .Z(N1607) );
  CAOR1X1 U19 ( .A(n12), .B(N1712), .C(N1483), .Z(N1603) );
  CAOR1X1 U20 ( .A(n12), .B(N1713), .C(N1483), .Z(N1599) );
  CAOR1X1 U21 ( .A(n12), .B(N1714), .C(N1483), .Z(N1595) );
  CAOR1X1 U22 ( .A(n12), .B(N1715), .C(N1483), .Z(N1591) );
  CAOR1X1 U23 ( .A(n12), .B(N1716), .C(N1483), .Z(N1587) );
  CAOR1X1 U24 ( .A(n12), .B(N1717), .C(N1483), .Z(N1583) );
  CAOR1X1 U25 ( .A(n12), .B(N1718), .C(N1483), .Z(N1579) );
  CAOR1X1 U26 ( .A(n12), .B(N1719), .C(N1483), .Z(N1575) );
  CAOR1X1 U27 ( .A(n12), .B(N1720), .C(N1483), .Z(N1571) );
  CAOR1X1 U28 ( .A(n12), .B(N1721), .C(N1483), .Z(N1567) );
  CAOR1X1 U29 ( .A(n12), .B(N1722), .C(N1483), .Z(N1563) );
  CAOR1X1 U30 ( .A(n12), .B(N1723), .C(N1483), .Z(N1559) );
  CAOR1X1 U31 ( .A(n12), .B(N1724), .C(N1483), .Z(N1555) );
  CAOR1X1 U32 ( .A(n12), .B(N1725), .C(N1483), .Z(N1551) );
  CAOR1X1 U33 ( .A(n12), .B(N1726), .C(N1483), .Z(N1547) );
  CAOR1X1 U34 ( .A(n12), .B(N1727), .C(N1483), .Z(N1543) );
  CAOR1X1 U35 ( .A(n12), .B(N1728), .C(N1483), .Z(N1539) );
  CAOR1X1 U36 ( .A(n12), .B(N1729), .C(N1483), .Z(N1535) );
  CAOR1X1 U37 ( .A(n12), .B(N1730), .C(N1483), .Z(N1531) );
  CAOR1X1 U38 ( .A(n12), .B(N1731), .C(N1483), .Z(N1527) );
  CAOR1X1 U39 ( .A(n12), .B(N1732), .C(N1483), .Z(N1523) );
  CNR2X1 U40 ( .A(n13), .B(n14), .Z(n12) );
  CAOR1X1 U42 ( .A(reset), .B(n652), .C(N1651), .Z(N1483) );
  CANR1XL U44 ( .A(n592), .B(N1037), .C(n14), .Z(N1482) );
  CND2X1 U49 ( .A(n19), .B(n20), .Z(N1351) );
  CND2X1 U50 ( .A(N249), .B(n13), .Z(n20) );
  CND2X1 U52 ( .A(n21), .B(n22), .Z(N1349) );
  CANR2X1 U54 ( .A(N119), .B(n652), .C(N592), .D(n18), .Z(n21) );
  CND2X1 U55 ( .A(n23), .B(n24), .Z(N1347) );
  CND2X1 U56 ( .A(N251), .B(n13), .Z(n24) );
  CND2X1 U58 ( .A(n25), .B(n26), .Z(N1345) );
  CND2X1 U61 ( .A(n27), .B(n28), .Z(N1343) );
  CND2X1 U62 ( .A(N253), .B(n13), .Z(n28) );
  CND2X1 U64 ( .A(n29), .B(n30), .Z(N1341) );
  CND2X1 U65 ( .A(N254), .B(n13), .Z(n30) );
  CANR2X1 U66 ( .A(N111), .B(n652), .C(N588), .D(n18), .Z(n29) );
  CND2X1 U67 ( .A(n31), .B(n32), .Z(N1339) );
  CND2X1 U68 ( .A(N255), .B(n13), .Z(n32) );
  CANR2X1 U69 ( .A(N109), .B(n652), .C(N587), .D(n18), .Z(n31) );
  CND2X1 U70 ( .A(n33), .B(n34), .Z(N1337) );
  CND2X1 U71 ( .A(N256), .B(n13), .Z(n34) );
  CANR2X1 U72 ( .A(N107), .B(n651), .C(N586), .D(n18), .Z(n33) );
  CND2X1 U73 ( .A(n35), .B(n36), .Z(N1335) );
  CND2X1 U74 ( .A(N257), .B(n13), .Z(n36) );
  CANR2X1 U75 ( .A(N105), .B(n651), .C(N585), .D(n18), .Z(n35) );
  CND2X1 U76 ( .A(n37), .B(n38), .Z(N1333) );
  CND2X1 U77 ( .A(N258), .B(n13), .Z(n38) );
  CANR2X1 U78 ( .A(N103), .B(n651), .C(N584), .D(n18), .Z(n37) );
  CND2X1 U79 ( .A(n39), .B(n40), .Z(N1331) );
  CND2X1 U80 ( .A(N259), .B(n13), .Z(n40) );
  CANR2X1 U81 ( .A(N101), .B(n651), .C(N583), .D(n18), .Z(n39) );
  CND2X1 U82 ( .A(n41), .B(n42), .Z(N1329) );
  CND2X1 U83 ( .A(N260), .B(n13), .Z(n42) );
  CANR2X1 U84 ( .A(N99), .B(n651), .C(N582), .D(n18), .Z(n41) );
  CND2X1 U85 ( .A(n43), .B(n44), .Z(N1327) );
  CND2X1 U86 ( .A(N261), .B(n13), .Z(n44) );
  CANR2X1 U87 ( .A(N97), .B(n651), .C(N581), .D(n18), .Z(n43) );
  CND2X1 U88 ( .A(n45), .B(n46), .Z(N1325) );
  CND2X1 U89 ( .A(N262), .B(n13), .Z(n46) );
  CANR2X1 U90 ( .A(N95), .B(n651), .C(N580), .D(n18), .Z(n45) );
  CND2X1 U91 ( .A(n47), .B(n48), .Z(N1323) );
  CND2X1 U92 ( .A(N263), .B(n13), .Z(n48) );
  CND2X1 U95 ( .A(N264), .B(n13), .Z(n50) );
  CND2X1 U97 ( .A(n51), .B(n52), .Z(N1319) );
  CND2X1 U98 ( .A(N265), .B(n13), .Z(n52) );
  CANR2X1 U99 ( .A(N89), .B(n651), .C(N577), .D(n18), .Z(n51) );
  CND2X1 U100 ( .A(n53), .B(n54), .Z(N1317) );
  CND2X1 U101 ( .A(N266), .B(n13), .Z(n54) );
  CND2X1 U104 ( .A(N267), .B(n13), .Z(n56) );
  CND2X1 U106 ( .A(n57), .B(n58), .Z(N1313) );
  CND2X1 U107 ( .A(N268), .B(n13), .Z(n58) );
  CANR2X1 U108 ( .A(N83), .B(n651), .C(N574), .D(n18), .Z(n57) );
  CND2X1 U109 ( .A(n59), .B(n60), .Z(N1311) );
  CND2X1 U110 ( .A(N269), .B(n13), .Z(n60) );
  CANR2X1 U111 ( .A(N81), .B(n651), .C(N573), .D(n18), .Z(n59) );
  CND2X1 U112 ( .A(n61), .B(n62), .Z(N1309) );
  CND2X1 U113 ( .A(N270), .B(n13), .Z(n62) );
  CANR2X1 U114 ( .A(N79), .B(n650), .C(N572), .D(n18), .Z(n61) );
  CND2X1 U115 ( .A(n63), .B(n64), .Z(N1307) );
  CND2X1 U116 ( .A(N271), .B(n13), .Z(n64) );
  CANR2X1 U117 ( .A(N77), .B(n650), .C(N571), .D(n18), .Z(n63) );
  CND2X1 U118 ( .A(n65), .B(n66), .Z(N1305) );
  CND2X1 U119 ( .A(N272), .B(n13), .Z(n66) );
  CANR2X1 U120 ( .A(N75), .B(n650), .C(N570), .D(n18), .Z(n65) );
  CND2X1 U121 ( .A(n67), .B(n68), .Z(N1303) );
  CND2X1 U122 ( .A(N273), .B(n13), .Z(n68) );
  CANR2X1 U123 ( .A(N73), .B(n650), .C(N569), .D(n18), .Z(n67) );
  CND2X1 U124 ( .A(n69), .B(n70), .Z(N1301) );
  CND2X1 U125 ( .A(N274), .B(n13), .Z(n70) );
  CANR2X1 U126 ( .A(N71), .B(n650), .C(N568), .D(n18), .Z(n69) );
  COND1XL U127 ( .A(n518), .B(N3), .C(n71), .Z(N1299) );
  COND1XL U129 ( .A(n518), .B(n552), .C(n72), .Z(N1297) );
  CANR2X1 U130 ( .A(N67), .B(n650), .C(N566), .D(n18), .Z(n72) );
  COND1XL U131 ( .A(n518), .B(N1688), .C(n73), .Z(N1295) );
  COND1XL U133 ( .A(n518), .B(N7), .C(n74), .Z(N1293) );
  COND1XL U135 ( .A(n518), .B(N6), .C(n75), .Z(N1291) );
  CAOR2X1 U138 ( .A(n78), .B(N1702), .C(\memory[31][2] ), .D(n77), .Z(N1283)
         );
  CAOR2X1 U141 ( .A(n80), .B(N1702), .C(\memory[31][0] ), .D(n77), .Z(N1279)
         );
  CND2X1 U142 ( .A(N1702), .B(n18), .Z(n77) );
  CIVX1 U143 ( .A(N1037), .Z(n18) );
  CND2X1 U144 ( .A(n81), .B(n82), .Z(N1277) );
  CND2X1 U145 ( .A(N711), .B(n650), .Z(n82) );
  CANR2X1 U146 ( .A(\memory[30][3] ), .B(n83), .C(n76), .D(N1703), .Z(n81) );
  CND2X1 U147 ( .A(n84), .B(n85), .Z(N1275) );
  CND2X1 U148 ( .A(N712), .B(n650), .Z(n85) );
  CANR2X1 U149 ( .A(\memory[30][2] ), .B(n83), .C(n78), .D(N1703), .Z(n84) );
  CND2X1 U150 ( .A(n86), .B(n87), .Z(N1273) );
  CND2X1 U151 ( .A(N713), .B(n650), .Z(n87) );
  CANR2X1 U152 ( .A(\memory[30][1] ), .B(n83), .C(n79), .D(N1703), .Z(n86) );
  CND2X1 U153 ( .A(n88), .B(n89), .Z(N1271) );
  CND2X1 U154 ( .A(N714), .B(n649), .Z(n89) );
  CANR2X1 U155 ( .A(\memory[30][0] ), .B(n83), .C(n80), .D(N1703), .Z(n88) );
  COND1XL U156 ( .A(N1703), .B(n90), .C(wr_enable), .Z(n83) );
  CND2X1 U157 ( .A(n91), .B(n92), .Z(N1269) );
  CND2X1 U158 ( .A(N707), .B(n649), .Z(n92) );
  CANR2X1 U159 ( .A(\memory[29][3] ), .B(n93), .C(n76), .D(N1704), .Z(n91) );
  CND2X1 U160 ( .A(n94), .B(n95), .Z(N1267) );
  CND2X1 U161 ( .A(N708), .B(n649), .Z(n95) );
  CANR2X1 U162 ( .A(\memory[29][2] ), .B(n93), .C(n78), .D(N1704), .Z(n94) );
  CND2X1 U163 ( .A(n96), .B(n97), .Z(N1265) );
  CND2X1 U164 ( .A(N709), .B(n649), .Z(n97) );
  CANR2X1 U165 ( .A(\memory[29][1] ), .B(n93), .C(n79), .D(N1704), .Z(n96) );
  CND2X1 U166 ( .A(n98), .B(n99), .Z(N1263) );
  CND2X1 U167 ( .A(N710), .B(n649), .Z(n99) );
  CANR2X1 U168 ( .A(\memory[29][0] ), .B(n93), .C(n80), .D(N1704), .Z(n98) );
  COND1XL U169 ( .A(N1704), .B(n90), .C(wr_enable), .Z(n93) );
  CND2X1 U170 ( .A(n100), .B(n101), .Z(N1261) );
  CND2X1 U171 ( .A(N703), .B(n649), .Z(n101) );
  CANR2X1 U172 ( .A(\memory[28][3] ), .B(n102), .C(n76), .D(N1705), .Z(n100)
         );
  CND2X1 U173 ( .A(n103), .B(n104), .Z(N1259) );
  CND2X1 U174 ( .A(N704), .B(n649), .Z(n104) );
  CANR2X1 U175 ( .A(\memory[28][2] ), .B(n102), .C(n78), .D(N1705), .Z(n103)
         );
  CND2X1 U176 ( .A(n105), .B(n106), .Z(N1257) );
  CND2X1 U177 ( .A(N705), .B(n649), .Z(n106) );
  CANR2X1 U178 ( .A(\memory[28][1] ), .B(n102), .C(n79), .D(N1705), .Z(n105)
         );
  CND2X1 U179 ( .A(n107), .B(n108), .Z(N1255) );
  CND2X1 U180 ( .A(N706), .B(n649), .Z(n108) );
  CANR2X1 U181 ( .A(\memory[28][0] ), .B(n102), .C(n80), .D(N1705), .Z(n107)
         );
  COND1XL U182 ( .A(N1705), .B(n90), .C(wr_enable), .Z(n102) );
  CND2X1 U183 ( .A(n109), .B(n110), .Z(N1253) );
  CND2X1 U184 ( .A(N699), .B(n649), .Z(n110) );
  CANR2X1 U185 ( .A(\memory[27][3] ), .B(n111), .C(n76), .D(N1706), .Z(n109)
         );
  CND2X1 U186 ( .A(n112), .B(n113), .Z(N1251) );
  CND2X1 U187 ( .A(N700), .B(n649), .Z(n113) );
  CANR2X1 U188 ( .A(\memory[27][2] ), .B(n111), .C(n78), .D(N1706), .Z(n112)
         );
  CND2X1 U189 ( .A(n114), .B(n115), .Z(N1249) );
  CND2X1 U190 ( .A(N701), .B(n649), .Z(n115) );
  CANR2X1 U191 ( .A(\memory[27][1] ), .B(n111), .C(n79), .D(N1706), .Z(n114)
         );
  CND2X1 U192 ( .A(n116), .B(n117), .Z(N1247) );
  CND2X1 U193 ( .A(N702), .B(n649), .Z(n117) );
  CANR2X1 U194 ( .A(\memory[27][0] ), .B(n111), .C(n80), .D(N1706), .Z(n116)
         );
  COND1XL U195 ( .A(N1706), .B(n90), .C(wr_enable), .Z(n111) );
  CND2X1 U196 ( .A(n118), .B(n119), .Z(N1245) );
  CND2X1 U197 ( .A(N695), .B(n648), .Z(n119) );
  CANR2X1 U198 ( .A(\memory[26][3] ), .B(n120), .C(n76), .D(N1707), .Z(n118)
         );
  CND2X1 U199 ( .A(n121), .B(n122), .Z(N1243) );
  CND2X1 U200 ( .A(N696), .B(n648), .Z(n122) );
  CANR2X1 U201 ( .A(\memory[26][2] ), .B(n120), .C(n78), .D(N1707), .Z(n121)
         );
  CND2X1 U202 ( .A(n123), .B(n124), .Z(N1241) );
  CND2X1 U203 ( .A(N697), .B(n648), .Z(n124) );
  CANR2X1 U204 ( .A(\memory[26][1] ), .B(n120), .C(n79), .D(N1707), .Z(n123)
         );
  CND2X1 U205 ( .A(n125), .B(n126), .Z(N1239) );
  CND2X1 U206 ( .A(N698), .B(n648), .Z(n126) );
  CANR2X1 U207 ( .A(\memory[26][0] ), .B(n120), .C(n80), .D(N1707), .Z(n125)
         );
  COND1XL U208 ( .A(N1707), .B(n90), .C(wr_enable), .Z(n120) );
  CND2X1 U209 ( .A(n127), .B(n128), .Z(N1237) );
  CND2X1 U210 ( .A(N691), .B(n648), .Z(n128) );
  CANR2X1 U211 ( .A(\memory[25][3] ), .B(n129), .C(n76), .D(N1708), .Z(n127)
         );
  CND2X1 U212 ( .A(n130), .B(n131), .Z(N1235) );
  CND2X1 U213 ( .A(N692), .B(n648), .Z(n131) );
  CANR2X1 U214 ( .A(\memory[25][2] ), .B(n129), .C(n78), .D(N1708), .Z(n130)
         );
  CND2X1 U215 ( .A(n132), .B(n133), .Z(N1233) );
  CND2X1 U216 ( .A(N693), .B(n648), .Z(n133) );
  CANR2X1 U217 ( .A(\memory[25][1] ), .B(n129), .C(n79), .D(N1708), .Z(n132)
         );
  CND2X1 U218 ( .A(n134), .B(n135), .Z(N1231) );
  CND2X1 U219 ( .A(N694), .B(n648), .Z(n135) );
  CANR2X1 U220 ( .A(\memory[25][0] ), .B(n129), .C(n80), .D(N1708), .Z(n134)
         );
  COND1XL U221 ( .A(N1708), .B(n90), .C(wr_enable), .Z(n129) );
  CND2X1 U222 ( .A(n136), .B(n137), .Z(N1229) );
  CND2X1 U223 ( .A(N687), .B(n648), .Z(n137) );
  CANR2X1 U224 ( .A(\memory[24][3] ), .B(n138), .C(n76), .D(N1709), .Z(n136)
         );
  CND2X1 U225 ( .A(n139), .B(n140), .Z(N1227) );
  CND2X1 U226 ( .A(N688), .B(n648), .Z(n140) );
  CANR2X1 U227 ( .A(\memory[24][2] ), .B(n138), .C(n78), .D(N1709), .Z(n139)
         );
  CND2X1 U228 ( .A(n141), .B(n142), .Z(N1225) );
  CND2X1 U229 ( .A(N689), .B(n648), .Z(n142) );
  CANR2X1 U230 ( .A(\memory[24][1] ), .B(n138), .C(n79), .D(N1709), .Z(n141)
         );
  CND2X1 U231 ( .A(n143), .B(n144), .Z(N1223) );
  CND2X1 U232 ( .A(N690), .B(n648), .Z(n144) );
  CANR2X1 U233 ( .A(\memory[24][0] ), .B(n138), .C(n80), .D(N1709), .Z(n143)
         );
  COND1XL U234 ( .A(N1709), .B(n90), .C(wr_enable), .Z(n138) );
  CND2X1 U235 ( .A(n145), .B(n146), .Z(N1221) );
  CND2X1 U236 ( .A(N683), .B(n648), .Z(n146) );
  CANR2X1 U237 ( .A(\memory[23][3] ), .B(n147), .C(n76), .D(N1710), .Z(n145)
         );
  CND2X1 U238 ( .A(n148), .B(n149), .Z(N1219) );
  CND2X1 U239 ( .A(N684), .B(n647), .Z(n149) );
  CANR2X1 U240 ( .A(\memory[23][2] ), .B(n147), .C(n78), .D(N1710), .Z(n148)
         );
  CND2X1 U241 ( .A(n150), .B(n151), .Z(N1217) );
  CND2X1 U242 ( .A(N685), .B(n647), .Z(n151) );
  CANR2X1 U243 ( .A(\memory[23][1] ), .B(n147), .C(n79), .D(N1710), .Z(n150)
         );
  CND2X1 U244 ( .A(n152), .B(n153), .Z(N1215) );
  CND2X1 U245 ( .A(N686), .B(n647), .Z(n153) );
  CANR2X1 U246 ( .A(\memory[23][0] ), .B(n147), .C(n80), .D(N1710), .Z(n152)
         );
  COND1XL U247 ( .A(N1710), .B(n90), .C(wr_enable), .Z(n147) );
  CND2X1 U248 ( .A(n154), .B(n155), .Z(N1213) );
  CND2X1 U249 ( .A(N679), .B(n647), .Z(n155) );
  CANR2X1 U250 ( .A(\memory[22][3] ), .B(n156), .C(n76), .D(N1711), .Z(n154)
         );
  CND2X1 U251 ( .A(n157), .B(n158), .Z(N1211) );
  CND2X1 U252 ( .A(N680), .B(n647), .Z(n158) );
  CANR2X1 U253 ( .A(\memory[22][2] ), .B(n156), .C(n78), .D(N1711), .Z(n157)
         );
  CND2X1 U254 ( .A(n159), .B(n160), .Z(N1209) );
  CND2X1 U255 ( .A(N681), .B(n647), .Z(n160) );
  CANR2X1 U256 ( .A(\memory[22][1] ), .B(n156), .C(n79), .D(N1711), .Z(n159)
         );
  CND2X1 U257 ( .A(n161), .B(n162), .Z(N1207) );
  CND2X1 U258 ( .A(N682), .B(n647), .Z(n162) );
  CANR2X1 U259 ( .A(\memory[22][0] ), .B(n156), .C(n80), .D(N1711), .Z(n161)
         );
  COND1XL U260 ( .A(N1711), .B(n90), .C(wr_enable), .Z(n156) );
  CND2X1 U261 ( .A(n163), .B(n164), .Z(N1205) );
  CND2X1 U262 ( .A(N675), .B(n647), .Z(n164) );
  CANR2X1 U263 ( .A(\memory[21][3] ), .B(n165), .C(n76), .D(N1712), .Z(n163)
         );
  CND2X1 U264 ( .A(n166), .B(n167), .Z(N1203) );
  CND2X1 U265 ( .A(N676), .B(n647), .Z(n167) );
  CANR2X1 U266 ( .A(\memory[21][2] ), .B(n165), .C(n78), .D(N1712), .Z(n166)
         );
  CND2X1 U267 ( .A(n168), .B(n169), .Z(N1201) );
  CND2X1 U268 ( .A(N677), .B(n647), .Z(n169) );
  CANR2X1 U269 ( .A(\memory[21][1] ), .B(n165), .C(n79), .D(N1712), .Z(n168)
         );
  CND2X1 U270 ( .A(n170), .B(n171), .Z(N1199) );
  CND2X1 U271 ( .A(N678), .B(n647), .Z(n171) );
  CANR2X1 U272 ( .A(\memory[21][0] ), .B(n165), .C(n80), .D(N1712), .Z(n170)
         );
  COND1XL U273 ( .A(N1712), .B(n90), .C(wr_enable), .Z(n165) );
  CND2X1 U274 ( .A(n172), .B(n173), .Z(N1197) );
  CND2X1 U275 ( .A(N671), .B(n647), .Z(n173) );
  CANR2X1 U276 ( .A(\memory[20][3] ), .B(n174), .C(n76), .D(N1713), .Z(n172)
         );
  CND2X1 U277 ( .A(n175), .B(n176), .Z(N1195) );
  CND2X1 U278 ( .A(N672), .B(n647), .Z(n176) );
  CANR2X1 U279 ( .A(\memory[20][2] ), .B(n174), .C(n78), .D(N1713), .Z(n175)
         );
  CND2X1 U280 ( .A(n177), .B(n178), .Z(N1193) );
  CND2X1 U281 ( .A(N673), .B(n646), .Z(n178) );
  CANR2X1 U282 ( .A(\memory[20][1] ), .B(n174), .C(n79), .D(N1713), .Z(n177)
         );
  CND2X1 U283 ( .A(n179), .B(n180), .Z(N1191) );
  CND2X1 U284 ( .A(N674), .B(n646), .Z(n180) );
  CANR2X1 U285 ( .A(\memory[20][0] ), .B(n174), .C(n80), .D(N1713), .Z(n179)
         );
  COND1XL U286 ( .A(N1713), .B(n90), .C(wr_enable), .Z(n174) );
  CND2X1 U287 ( .A(n181), .B(n182), .Z(N1189) );
  CND2X1 U288 ( .A(N667), .B(n646), .Z(n182) );
  CANR2X1 U289 ( .A(\memory[19][3] ), .B(n183), .C(n76), .D(N1714), .Z(n181)
         );
  CND2X1 U290 ( .A(n184), .B(n185), .Z(N1187) );
  CND2X1 U291 ( .A(N668), .B(n646), .Z(n185) );
  CANR2X1 U292 ( .A(\memory[19][2] ), .B(n183), .C(n78), .D(N1714), .Z(n184)
         );
  CND2X1 U293 ( .A(n186), .B(n187), .Z(N1185) );
  CND2X1 U294 ( .A(N669), .B(n646), .Z(n187) );
  CANR2X1 U295 ( .A(\memory[19][1] ), .B(n183), .C(n79), .D(N1714), .Z(n186)
         );
  CND2X1 U296 ( .A(n188), .B(n189), .Z(N1183) );
  CND2X1 U297 ( .A(N670), .B(n646), .Z(n189) );
  CANR2X1 U298 ( .A(\memory[19][0] ), .B(n183), .C(n80), .D(N1714), .Z(n188)
         );
  COND1XL U299 ( .A(N1714), .B(n90), .C(wr_enable), .Z(n183) );
  CND2X1 U300 ( .A(n190), .B(n191), .Z(N1181) );
  CND2X1 U301 ( .A(N663), .B(n646), .Z(n191) );
  CANR2X1 U302 ( .A(\memory[18][3] ), .B(n192), .C(n76), .D(N1715), .Z(n190)
         );
  CND2X1 U303 ( .A(n193), .B(n194), .Z(N1179) );
  CND2X1 U304 ( .A(N664), .B(n646), .Z(n194) );
  CANR2X1 U305 ( .A(\memory[18][2] ), .B(n192), .C(n78), .D(N1715), .Z(n193)
         );
  CND2X1 U306 ( .A(n195), .B(n196), .Z(N1177) );
  CND2X1 U307 ( .A(N665), .B(n646), .Z(n196) );
  CANR2X1 U308 ( .A(\memory[18][1] ), .B(n192), .C(n79), .D(N1715), .Z(n195)
         );
  CND2X1 U309 ( .A(n197), .B(n198), .Z(N1175) );
  CND2X1 U310 ( .A(N666), .B(n646), .Z(n198) );
  CANR2X1 U311 ( .A(\memory[18][0] ), .B(n192), .C(n80), .D(N1715), .Z(n197)
         );
  COND1XL U312 ( .A(N1715), .B(n90), .C(wr_enable), .Z(n192) );
  CND2X1 U313 ( .A(n199), .B(n200), .Z(N1173) );
  CND2X1 U314 ( .A(N659), .B(n646), .Z(n200) );
  CANR2X1 U315 ( .A(\memory[17][3] ), .B(n201), .C(n76), .D(N1716), .Z(n199)
         );
  CND2X1 U316 ( .A(n202), .B(n203), .Z(N1171) );
  CND2X1 U317 ( .A(N660), .B(n646), .Z(n203) );
  CANR2X1 U318 ( .A(\memory[17][2] ), .B(n201), .C(n78), .D(N1716), .Z(n202)
         );
  CND2X1 U319 ( .A(n204), .B(n205), .Z(N1169) );
  CND2X1 U320 ( .A(N661), .B(n646), .Z(n205) );
  CANR2X1 U321 ( .A(\memory[17][1] ), .B(n201), .C(n79), .D(N1716), .Z(n204)
         );
  CND2X1 U322 ( .A(n206), .B(n207), .Z(N1167) );
  CND2X1 U323 ( .A(N662), .B(n645), .Z(n207) );
  CANR2X1 U324 ( .A(\memory[17][0] ), .B(n201), .C(n80), .D(N1716), .Z(n206)
         );
  COND1XL U325 ( .A(N1716), .B(n90), .C(wr_enable), .Z(n201) );
  CND2X1 U326 ( .A(n208), .B(n209), .Z(N1165) );
  CND2X1 U327 ( .A(N655), .B(n645), .Z(n209) );
  CANR2X1 U328 ( .A(\memory[16][3] ), .B(n210), .C(n76), .D(N1717), .Z(n208)
         );
  CND2X1 U329 ( .A(n211), .B(n212), .Z(N1163) );
  CND2X1 U330 ( .A(N656), .B(n645), .Z(n212) );
  CANR2X1 U331 ( .A(\memory[16][2] ), .B(n210), .C(n78), .D(N1717), .Z(n211)
         );
  CND2X1 U332 ( .A(n213), .B(n214), .Z(N1161) );
  CND2X1 U333 ( .A(N657), .B(n645), .Z(n214) );
  CANR2X1 U334 ( .A(\memory[16][1] ), .B(n210), .C(n79), .D(N1717), .Z(n213)
         );
  CND2X1 U335 ( .A(n215), .B(n216), .Z(N1159) );
  CND2X1 U336 ( .A(N658), .B(n645), .Z(n216) );
  CANR2X1 U337 ( .A(\memory[16][0] ), .B(n210), .C(n80), .D(N1717), .Z(n215)
         );
  COND1XL U338 ( .A(N1717), .B(n90), .C(wr_enable), .Z(n210) );
  CND2X1 U339 ( .A(n217), .B(n218), .Z(N1157) );
  CND2X1 U340 ( .A(N651), .B(n645), .Z(n218) );
  CANR2X1 U341 ( .A(\memory[15][3] ), .B(n219), .C(n76), .D(N1718), .Z(n217)
         );
  CND2X1 U342 ( .A(n220), .B(n221), .Z(N1155) );
  CND2X1 U343 ( .A(N652), .B(n645), .Z(n221) );
  CANR2X1 U344 ( .A(\memory[15][2] ), .B(n219), .C(n78), .D(N1718), .Z(n220)
         );
  CND2X1 U345 ( .A(n222), .B(n223), .Z(N1153) );
  CND2X1 U346 ( .A(N653), .B(n645), .Z(n223) );
  CANR2X1 U347 ( .A(\memory[15][1] ), .B(n219), .C(n79), .D(N1718), .Z(n222)
         );
  CND2X1 U348 ( .A(n224), .B(n225), .Z(N1151) );
  CND2X1 U349 ( .A(N654), .B(n645), .Z(n225) );
  CANR2X1 U350 ( .A(\memory[15][0] ), .B(n219), .C(n80), .D(N1718), .Z(n224)
         );
  COND1XL U351 ( .A(N1718), .B(n90), .C(wr_enable), .Z(n219) );
  CND2X1 U352 ( .A(n226), .B(n227), .Z(N1149) );
  CND2X1 U353 ( .A(N647), .B(n645), .Z(n227) );
  CANR2X1 U354 ( .A(\memory[14][3] ), .B(n228), .C(n76), .D(N1719), .Z(n226)
         );
  CND2X1 U355 ( .A(n229), .B(n230), .Z(N1147) );
  CND2X1 U356 ( .A(N648), .B(n645), .Z(n230) );
  CANR2X1 U357 ( .A(\memory[14][2] ), .B(n228), .C(n78), .D(N1719), .Z(n229)
         );
  CND2X1 U358 ( .A(n231), .B(n232), .Z(N1145) );
  CND2X1 U359 ( .A(N649), .B(n645), .Z(n232) );
  CANR2X1 U360 ( .A(\memory[14][1] ), .B(n228), .C(n79), .D(N1719), .Z(n231)
         );
  CND2X1 U361 ( .A(n233), .B(n234), .Z(N1143) );
  CND2X1 U362 ( .A(N650), .B(n645), .Z(n234) );
  CANR2X1 U363 ( .A(\memory[14][0] ), .B(n228), .C(n80), .D(N1719), .Z(n233)
         );
  COND1XL U364 ( .A(N1719), .B(n90), .C(wr_enable), .Z(n228) );
  CND2X1 U365 ( .A(n235), .B(n236), .Z(N1141) );
  CND2X1 U366 ( .A(N643), .B(n644), .Z(n236) );
  CANR2X1 U367 ( .A(\memory[13][3] ), .B(n237), .C(n76), .D(N1720), .Z(n235)
         );
  CND2X1 U368 ( .A(n238), .B(n239), .Z(N1139) );
  CND2X1 U369 ( .A(N644), .B(n644), .Z(n239) );
  CANR2X1 U370 ( .A(\memory[13][2] ), .B(n237), .C(n78), .D(N1720), .Z(n238)
         );
  CND2X1 U371 ( .A(n240), .B(n241), .Z(N1137) );
  CND2X1 U372 ( .A(N645), .B(n644), .Z(n241) );
  CANR2X1 U373 ( .A(\memory[13][1] ), .B(n237), .C(n79), .D(N1720), .Z(n240)
         );
  CND2X1 U374 ( .A(n242), .B(n243), .Z(N1135) );
  CND2X1 U375 ( .A(N646), .B(n644), .Z(n243) );
  CANR2X1 U376 ( .A(\memory[13][0] ), .B(n237), .C(n80), .D(N1720), .Z(n242)
         );
  COND1XL U377 ( .A(N1720), .B(n90), .C(wr_enable), .Z(n237) );
  CND2X1 U378 ( .A(n244), .B(n245), .Z(N1133) );
  CND2X1 U379 ( .A(N639), .B(n644), .Z(n245) );
  CANR2X1 U380 ( .A(\memory[12][3] ), .B(n246), .C(n76), .D(N1721), .Z(n244)
         );
  CND2X1 U381 ( .A(n247), .B(n248), .Z(N1131) );
  CND2X1 U382 ( .A(N640), .B(n644), .Z(n248) );
  CANR2X1 U383 ( .A(\memory[12][2] ), .B(n246), .C(n78), .D(N1721), .Z(n247)
         );
  CND2X1 U384 ( .A(n249), .B(n250), .Z(N1129) );
  CND2X1 U385 ( .A(N641), .B(n644), .Z(n250) );
  CANR2X1 U386 ( .A(\memory[12][1] ), .B(n246), .C(n79), .D(N1721), .Z(n249)
         );
  CND2X1 U387 ( .A(n251), .B(n252), .Z(N1127) );
  CND2X1 U388 ( .A(N642), .B(n644), .Z(n252) );
  CANR2X1 U389 ( .A(\memory[12][0] ), .B(n246), .C(n80), .D(N1721), .Z(n251)
         );
  COND1XL U390 ( .A(N1721), .B(n90), .C(wr_enable), .Z(n246) );
  CND2X1 U391 ( .A(n253), .B(n254), .Z(N1125) );
  CND2X1 U392 ( .A(N635), .B(n644), .Z(n254) );
  CANR2X1 U393 ( .A(\memory[11][3] ), .B(n255), .C(n76), .D(N1722), .Z(n253)
         );
  CND2X1 U394 ( .A(n256), .B(n257), .Z(N1123) );
  CND2X1 U395 ( .A(N636), .B(n644), .Z(n257) );
  CANR2X1 U396 ( .A(\memory[11][2] ), .B(n255), .C(n78), .D(N1722), .Z(n256)
         );
  CND2X1 U397 ( .A(n258), .B(n259), .Z(N1121) );
  CND2X1 U398 ( .A(N637), .B(n644), .Z(n259) );
  CANR2X1 U399 ( .A(\memory[11][1] ), .B(n255), .C(n79), .D(N1722), .Z(n258)
         );
  CND2X1 U400 ( .A(n260), .B(n261), .Z(N1119) );
  CND2X1 U401 ( .A(N638), .B(n644), .Z(n261) );
  CANR2X1 U402 ( .A(\memory[11][0] ), .B(n255), .C(n80), .D(N1722), .Z(n260)
         );
  COND1XL U403 ( .A(N1722), .B(n90), .C(wr_enable), .Z(n255) );
  CND2X1 U404 ( .A(n262), .B(n263), .Z(N1117) );
  CND2X1 U405 ( .A(N631), .B(n644), .Z(n263) );
  CANR2X1 U406 ( .A(\memory[10][3] ), .B(n264), .C(n76), .D(N1723), .Z(n262)
         );
  CND2X1 U407 ( .A(n265), .B(n266), .Z(N1115) );
  CND2X1 U408 ( .A(N632), .B(n643), .Z(n266) );
  CANR2X1 U409 ( .A(\memory[10][2] ), .B(n264), .C(n78), .D(N1723), .Z(n265)
         );
  CND2X1 U410 ( .A(n267), .B(n268), .Z(N1113) );
  CND2X1 U411 ( .A(N633), .B(n643), .Z(n268) );
  CANR2X1 U412 ( .A(\memory[10][1] ), .B(n264), .C(n79), .D(N1723), .Z(n267)
         );
  CND2X1 U413 ( .A(n269), .B(n270), .Z(N1111) );
  CND2X1 U414 ( .A(N634), .B(n643), .Z(n270) );
  CANR2X1 U415 ( .A(\memory[10][0] ), .B(n264), .C(n80), .D(N1723), .Z(n269)
         );
  COND1XL U416 ( .A(N1723), .B(n90), .C(wr_enable), .Z(n264) );
  CND2X1 U417 ( .A(n271), .B(n272), .Z(N1109) );
  CND2X1 U418 ( .A(N627), .B(n643), .Z(n272) );
  CANR2X1 U419 ( .A(\memory[9][3] ), .B(n273), .C(n76), .D(N1724), .Z(n271) );
  CND2X1 U420 ( .A(n274), .B(n275), .Z(N1107) );
  CND2X1 U421 ( .A(N628), .B(n643), .Z(n275) );
  CANR2X1 U422 ( .A(\memory[9][2] ), .B(n273), .C(n78), .D(N1724), .Z(n274) );
  CND2X1 U423 ( .A(n276), .B(n277), .Z(N1105) );
  CND2X1 U424 ( .A(N629), .B(n643), .Z(n277) );
  CANR2X1 U425 ( .A(\memory[9][1] ), .B(n273), .C(n79), .D(N1724), .Z(n276) );
  CND2X1 U426 ( .A(n278), .B(n279), .Z(N1103) );
  CND2X1 U427 ( .A(N630), .B(n643), .Z(n279) );
  CANR2X1 U428 ( .A(\memory[9][0] ), .B(n273), .C(n80), .D(N1724), .Z(n278) );
  COND1XL U429 ( .A(N1724), .B(n90), .C(wr_enable), .Z(n273) );
  CND2X1 U430 ( .A(n280), .B(n281), .Z(N1101) );
  CND2X1 U431 ( .A(N623), .B(n643), .Z(n281) );
  CANR2X1 U432 ( .A(\memory[8][3] ), .B(n282), .C(n76), .D(N1725), .Z(n280) );
  CND2X1 U433 ( .A(n283), .B(n284), .Z(N1099) );
  CND2X1 U434 ( .A(N624), .B(n643), .Z(n284) );
  CANR2X1 U435 ( .A(\memory[8][2] ), .B(n282), .C(n78), .D(N1725), .Z(n283) );
  CND2X1 U436 ( .A(n285), .B(n286), .Z(N1097) );
  CND2X1 U437 ( .A(N625), .B(n643), .Z(n286) );
  CANR2X1 U438 ( .A(\memory[8][1] ), .B(n282), .C(n79), .D(N1725), .Z(n285) );
  CND2X1 U439 ( .A(n287), .B(n288), .Z(N1095) );
  CND2X1 U440 ( .A(N626), .B(n643), .Z(n288) );
  CANR2X1 U441 ( .A(\memory[8][0] ), .B(n282), .C(n80), .D(N1725), .Z(n287) );
  COND1XL U442 ( .A(N1725), .B(n90), .C(wr_enable), .Z(n282) );
  CND2X1 U443 ( .A(n289), .B(n290), .Z(N1093) );
  CND2X1 U444 ( .A(N619), .B(n643), .Z(n290) );
  CANR2X1 U445 ( .A(\memory[7][3] ), .B(n291), .C(n76), .D(N1726), .Z(n289) );
  CND2X1 U446 ( .A(n292), .B(n293), .Z(N1091) );
  CND2X1 U447 ( .A(N620), .B(n643), .Z(n293) );
  CANR2X1 U448 ( .A(\memory[7][2] ), .B(n291), .C(n78), .D(N1726), .Z(n292) );
  CND2X1 U449 ( .A(n294), .B(n295), .Z(N1089) );
  CND2X1 U450 ( .A(N621), .B(n642), .Z(n295) );
  CANR2X1 U451 ( .A(\memory[7][1] ), .B(n291), .C(n79), .D(N1726), .Z(n294) );
  CND2X1 U452 ( .A(n296), .B(n297), .Z(N1087) );
  CND2X1 U453 ( .A(N622), .B(n642), .Z(n297) );
  CANR2X1 U454 ( .A(\memory[7][0] ), .B(n291), .C(n80), .D(N1726), .Z(n296) );
  COND1XL U455 ( .A(N1726), .B(n90), .C(wr_enable), .Z(n291) );
  CND2X1 U456 ( .A(n298), .B(n299), .Z(N1085) );
  CND2X1 U457 ( .A(N615), .B(n642), .Z(n299) );
  CANR2X1 U458 ( .A(\memory[6][3] ), .B(n300), .C(n76), .D(N1727), .Z(n298) );
  CND2X1 U459 ( .A(n301), .B(n302), .Z(N1083) );
  CND2X1 U460 ( .A(N616), .B(n642), .Z(n302) );
  CANR2X1 U461 ( .A(\memory[6][2] ), .B(n300), .C(n78), .D(N1727), .Z(n301) );
  CND2X1 U462 ( .A(n303), .B(n304), .Z(N1081) );
  CND2X1 U463 ( .A(N617), .B(n642), .Z(n304) );
  CANR2X1 U464 ( .A(\memory[6][1] ), .B(n300), .C(n79), .D(N1727), .Z(n303) );
  CND2X1 U465 ( .A(n305), .B(n306), .Z(N1079) );
  CND2X1 U466 ( .A(N618), .B(n642), .Z(n306) );
  CANR2X1 U467 ( .A(\memory[6][0] ), .B(n300), .C(n80), .D(N1727), .Z(n305) );
  COND1XL U468 ( .A(N1727), .B(n90), .C(wr_enable), .Z(n300) );
  CND2X1 U469 ( .A(n307), .B(n308), .Z(N1077) );
  CND2X1 U470 ( .A(N611), .B(n642), .Z(n308) );
  CANR2X1 U471 ( .A(\memory[5][3] ), .B(n309), .C(n76), .D(N1728), .Z(n307) );
  CND2X1 U472 ( .A(n310), .B(n311), .Z(N1075) );
  CND2X1 U473 ( .A(N612), .B(n642), .Z(n311) );
  CANR2X1 U474 ( .A(\memory[5][2] ), .B(n309), .C(n78), .D(N1728), .Z(n310) );
  CND2X1 U475 ( .A(n312), .B(n313), .Z(N1073) );
  CND2X1 U476 ( .A(N613), .B(n642), .Z(n313) );
  CANR2X1 U477 ( .A(\memory[5][1] ), .B(n309), .C(n79), .D(N1728), .Z(n312) );
  CND2X1 U478 ( .A(n314), .B(n315), .Z(N1071) );
  CND2X1 U479 ( .A(N614), .B(n642), .Z(n315) );
  CANR2X1 U480 ( .A(\memory[5][0] ), .B(n309), .C(n80), .D(N1728), .Z(n314) );
  COND1XL U481 ( .A(N1728), .B(n90), .C(wr_enable), .Z(n309) );
  CND2X1 U482 ( .A(n316), .B(n317), .Z(N1069) );
  CND2X1 U483 ( .A(N607), .B(n642), .Z(n317) );
  CANR2X1 U484 ( .A(\memory[4][3] ), .B(n318), .C(n76), .D(N1729), .Z(n316) );
  CND2X1 U485 ( .A(n319), .B(n320), .Z(N1067) );
  CND2X1 U486 ( .A(N608), .B(n642), .Z(n320) );
  CANR2X1 U487 ( .A(\memory[4][2] ), .B(n318), .C(n78), .D(N1729), .Z(n319) );
  CND2X1 U488 ( .A(n321), .B(n322), .Z(N1065) );
  CND2X1 U489 ( .A(N609), .B(n642), .Z(n322) );
  CANR2X1 U490 ( .A(\memory[4][1] ), .B(n318), .C(n79), .D(N1729), .Z(n321) );
  CND2X1 U491 ( .A(n323), .B(n324), .Z(N1063) );
  CND2X1 U492 ( .A(N610), .B(n641), .Z(n324) );
  CANR2X1 U493 ( .A(\memory[4][0] ), .B(n318), .C(n80), .D(N1729), .Z(n323) );
  COND1XL U494 ( .A(N1729), .B(n90), .C(wr_enable), .Z(n318) );
  CND2X1 U495 ( .A(n325), .B(n326), .Z(N1061) );
  CND2X1 U496 ( .A(N603), .B(n641), .Z(n326) );
  CANR2X1 U497 ( .A(\memory[3][3] ), .B(n327), .C(n76), .D(N1730), .Z(n325) );
  CND2X1 U498 ( .A(n328), .B(n329), .Z(N1059) );
  CND2X1 U499 ( .A(N604), .B(n641), .Z(n329) );
  CANR2X1 U500 ( .A(\memory[3][2] ), .B(n327), .C(n78), .D(N1730), .Z(n328) );
  CND2X1 U501 ( .A(n330), .B(n331), .Z(N1057) );
  CND2X1 U502 ( .A(N605), .B(n641), .Z(n331) );
  CANR2X1 U503 ( .A(\memory[3][1] ), .B(n327), .C(n79), .D(N1730), .Z(n330) );
  CND2X1 U504 ( .A(n332), .B(n333), .Z(N1055) );
  CND2X1 U505 ( .A(N606), .B(n641), .Z(n333) );
  CANR2X1 U506 ( .A(\memory[3][0] ), .B(n327), .C(n80), .D(N1730), .Z(n332) );
  COND1XL U507 ( .A(N1730), .B(n90), .C(wr_enable), .Z(n327) );
  CND2X1 U508 ( .A(n334), .B(n335), .Z(N1053) );
  CND2X1 U509 ( .A(N599), .B(n641), .Z(n335) );
  CANR2X1 U510 ( .A(\memory[2][3] ), .B(n336), .C(n76), .D(N1731), .Z(n334) );
  CND2X1 U511 ( .A(n337), .B(n338), .Z(N1051) );
  CND2X1 U512 ( .A(N600), .B(n641), .Z(n338) );
  CANR2X1 U513 ( .A(\memory[2][2] ), .B(n336), .C(n78), .D(N1731), .Z(n337) );
  CND2X1 U514 ( .A(n339), .B(n340), .Z(N1049) );
  CND2X1 U515 ( .A(N601), .B(n641), .Z(n340) );
  CANR2X1 U516 ( .A(\memory[2][1] ), .B(n336), .C(n79), .D(N1731), .Z(n339) );
  CND2X1 U517 ( .A(n341), .B(n342), .Z(N1047) );
  CND2X1 U518 ( .A(N602), .B(n641), .Z(n342) );
  CANR2X1 U519 ( .A(\memory[2][0] ), .B(n336), .C(n80), .D(N1731), .Z(n341) );
  COND1XL U520 ( .A(N1731), .B(n90), .C(wr_enable), .Z(n336) );
  CND2X1 U521 ( .A(n343), .B(n344), .Z(N1045) );
  CND2X1 U522 ( .A(N595), .B(n641), .Z(n344) );
  CANR2X1 U523 ( .A(\memory[1][3] ), .B(n345), .C(n76), .D(N1732), .Z(n343) );
  CNR2IX1 U524 ( .B(data[3]), .A(N1037), .Z(n76) );
  CND2X1 U525 ( .A(n346), .B(n347), .Z(N1043) );
  CND2X1 U526 ( .A(N596), .B(n641), .Z(n347) );
  CANR2X1 U527 ( .A(\memory[1][2] ), .B(n345), .C(n78), .D(N1732), .Z(n346) );
  CND2X1 U529 ( .A(n348), .B(n349), .Z(N1041) );
  CND2X1 U530 ( .A(N597), .B(n641), .Z(n349) );
  CANR2X1 U531 ( .A(\memory[1][1] ), .B(n345), .C(n79), .D(N1732), .Z(n348) );
  CNR2IX1 U532 ( .B(data[1]), .A(N1037), .Z(n79) );
  CND2X1 U533 ( .A(n350), .B(n351), .Z(N1039) );
  CND2X1 U534 ( .A(N598), .B(n641), .Z(n351) );
  CANR2X1 U535 ( .A(\memory[1][0] ), .B(n345), .C(n80), .D(N1732), .Z(n350) );
  COND1XL U537 ( .A(N1732), .B(n90), .C(wr_enable), .Z(n345) );
  CIVX1 U538 ( .A(N282), .Z(n90) );
  CNR2X1 U540 ( .A(n13), .B(N282), .Z(N1035) );
  CIVX1 U541 ( .A(wr_enable), .Z(n13) );
  CMX2X1 U546 ( .A0(counter[1]), .A1(N1293), .S(N1519), .Z(n515) );
  CMX2X1 U547 ( .A0(counter[2]), .A1(N1295), .S(N1519), .Z(n514) );
  CMX2X1 U548 ( .A0(counter[3]), .A1(N1297), .S(N1519), .Z(n513) );
  CMX2X1 U549 ( .A0(counter[4]), .A1(N1299), .S(N1519), .Z(n512) );
  CMX2X1 U550 ( .A0(counter[5]), .A1(N1301), .S(N1519), .Z(n511) );
  CMX2X1 U552 ( .A0(counter[7]), .A1(N1305), .S(N1519), .Z(n509) );
  CMX2X1 U553 ( .A0(counter[8]), .A1(N1307), .S(N1519), .Z(n508) );
  CMX2X1 U554 ( .A0(counter[9]), .A1(N1309), .S(N1519), .Z(n507) );
  CMX2X1 U555 ( .A0(counter[10]), .A1(N1311), .S(N1519), .Z(n506) );
  CMX2X1 U556 ( .A0(counter[11]), .A1(N1313), .S(N1519), .Z(n505) );
  CMX2X1 U557 ( .A0(counter[12]), .A1(N1315), .S(N1519), .Z(n504) );
  CMX2X1 U558 ( .A0(counter[13]), .A1(N1317), .S(N1519), .Z(n503) );
  CMX2X1 U559 ( .A0(counter[14]), .A1(N1319), .S(N1519), .Z(n502) );
  CMX2X1 U560 ( .A0(counter[15]), .A1(N1321), .S(N1519), .Z(n501) );
  CMX2X1 U561 ( .A0(counter[16]), .A1(N1323), .S(N1519), .Z(n500) );
  CMX2X1 U562 ( .A0(counter[17]), .A1(N1325), .S(N1519), .Z(n499) );
  CMX2X1 U564 ( .A0(counter[19]), .A1(N1329), .S(N1519), .Z(n497) );
  CMX2X1 U565 ( .A0(counter[20]), .A1(N1331), .S(N1519), .Z(n496) );
  CMX2X1 U566 ( .A0(counter[21]), .A1(N1333), .S(N1519), .Z(n495) );
  CMX2X1 U572 ( .A0(counter[27]), .A1(N1345), .S(N1519), .Z(n489) );
  CMX2X1 U573 ( .A0(counter[28]), .A1(N1347), .S(N1519), .Z(n488) );
  CMX2X1 U580 ( .A0(\memory[0][0] ), .A1(N1039), .S(N1523), .Z(n481) );
  CMX2X1 U581 ( .A0(code[0]), .A1(\memory[0][0] ), .S(N1651), .Z(n480) );
  CMX2X1 U582 ( .A0(n519), .A1(N1041), .S(N1523), .Z(n479) );
  CMX2X1 U583 ( .A0(code[1]), .A1(n519), .S(N1651), .Z(n478) );
  CMX2X1 U584 ( .A0(\memory[0][2] ), .A1(N1043), .S(N1523), .Z(n477) );
  CMX2X1 U585 ( .A0(code[2]), .A1(\memory[0][2] ), .S(N1651), .Z(n476) );
  CMX2X1 U586 ( .A0(\memory[0][3] ), .A1(N1045), .S(N1523), .Z(n475) );
  CMX2X1 U587 ( .A0(code[3]), .A1(\memory[0][3] ), .S(N1651), .Z(n474) );
  CMX2X1 U588 ( .A0(\memory[1][0] ), .A1(N1047), .S(N1527), .Z(n473) );
  CMX2X1 U589 ( .A0(\memory[1][1] ), .A1(N1049), .S(N1527), .Z(n472) );
  CMX2X1 U590 ( .A0(\memory[1][2] ), .A1(N1051), .S(N1527), .Z(n471) );
  CMX2X1 U591 ( .A0(\memory[1][3] ), .A1(N1053), .S(N1527), .Z(n470) );
  CMX2X1 U592 ( .A0(\memory[2][0] ), .A1(N1055), .S(N1531), .Z(n469) );
  CMX2X1 U593 ( .A0(\memory[2][1] ), .A1(N1057), .S(N1531), .Z(n468) );
  CMX2X1 U594 ( .A0(\memory[2][2] ), .A1(N1059), .S(N1531), .Z(n467) );
  CMX2X1 U595 ( .A0(\memory[2][3] ), .A1(N1061), .S(N1531), .Z(n466) );
  CMX2X1 U596 ( .A0(\memory[3][0] ), .A1(N1063), .S(N1535), .Z(n465) );
  CMX2X1 U597 ( .A0(\memory[3][1] ), .A1(N1065), .S(N1535), .Z(n464) );
  CMX2X1 U598 ( .A0(\memory[3][2] ), .A1(N1067), .S(N1535), .Z(n463) );
  CMX2X1 U599 ( .A0(\memory[3][3] ), .A1(N1069), .S(N1535), .Z(n462) );
  CMX2X1 U600 ( .A0(\memory[4][0] ), .A1(N1071), .S(N1539), .Z(n461) );
  CMX2X1 U601 ( .A0(\memory[4][1] ), .A1(N1073), .S(N1539), .Z(n460) );
  CMX2X1 U602 ( .A0(\memory[4][2] ), .A1(N1075), .S(N1539), .Z(n459) );
  CMX2X1 U603 ( .A0(\memory[4][3] ), .A1(N1077), .S(N1539), .Z(n458) );
  CMX2X1 U604 ( .A0(\memory[5][0] ), .A1(N1079), .S(N1543), .Z(n457) );
  CMX2X1 U605 ( .A0(\memory[5][1] ), .A1(N1081), .S(N1543), .Z(n456) );
  CMX2X1 U606 ( .A0(\memory[5][2] ), .A1(N1083), .S(N1543), .Z(n455) );
  CMX2X1 U607 ( .A0(\memory[5][3] ), .A1(N1085), .S(N1543), .Z(n454) );
  CMX2X1 U608 ( .A0(\memory[6][0] ), .A1(N1087), .S(N1547), .Z(n453) );
  CMX2X1 U609 ( .A0(\memory[6][1] ), .A1(N1089), .S(N1547), .Z(n452) );
  CMX2X1 U610 ( .A0(\memory[6][2] ), .A1(N1091), .S(N1547), .Z(n451) );
  CMX2X1 U611 ( .A0(\memory[6][3] ), .A1(N1093), .S(N1547), .Z(n450) );
  CMX2X1 U612 ( .A0(\memory[7][0] ), .A1(N1095), .S(N1551), .Z(n449) );
  CMX2X1 U613 ( .A0(\memory[7][1] ), .A1(N1097), .S(N1551), .Z(n448) );
  CMX2X1 U614 ( .A0(\memory[7][2] ), .A1(N1099), .S(N1551), .Z(n447) );
  CMX2X1 U615 ( .A0(\memory[7][3] ), .A1(N1101), .S(N1551), .Z(n446) );
  CMX2X1 U616 ( .A0(\memory[8][0] ), .A1(N1103), .S(N1555), .Z(n445) );
  CMX2X1 U617 ( .A0(\memory[8][1] ), .A1(N1105), .S(N1555), .Z(n444) );
  CMX2X1 U618 ( .A0(\memory[8][2] ), .A1(N1107), .S(N1555), .Z(n443) );
  CMX2X1 U619 ( .A0(\memory[8][3] ), .A1(N1109), .S(N1555), .Z(n442) );
  CMX2X1 U620 ( .A0(\memory[9][0] ), .A1(N1111), .S(N1559), .Z(n441) );
  CMX2X1 U621 ( .A0(\memory[9][1] ), .A1(N1113), .S(N1559), .Z(n440) );
  CMX2X1 U622 ( .A0(\memory[9][2] ), .A1(N1115), .S(N1559), .Z(n439) );
  CMX2X1 U623 ( .A0(\memory[9][3] ), .A1(N1117), .S(N1559), .Z(n438) );
  CMX2X1 U624 ( .A0(\memory[10][0] ), .A1(N1119), .S(N1563), .Z(n437) );
  CMX2X1 U625 ( .A0(\memory[10][1] ), .A1(N1121), .S(N1563), .Z(n436) );
  CMX2X1 U626 ( .A0(\memory[10][2] ), .A1(N1123), .S(N1563), .Z(n435) );
  CMX2X1 U627 ( .A0(\memory[10][3] ), .A1(N1125), .S(N1563), .Z(n434) );
  CMX2X1 U628 ( .A0(\memory[11][0] ), .A1(N1127), .S(N1567), .Z(n433) );
  CMX2X1 U629 ( .A0(\memory[11][1] ), .A1(N1129), .S(N1567), .Z(n432) );
  CMX2X1 U630 ( .A0(\memory[11][2] ), .A1(N1131), .S(N1567), .Z(n431) );
  CMX2X1 U631 ( .A0(\memory[11][3] ), .A1(N1133), .S(N1567), .Z(n430) );
  CMX2X1 U632 ( .A0(\memory[12][0] ), .A1(N1135), .S(N1571), .Z(n429) );
  CMX2X1 U633 ( .A0(\memory[12][1] ), .A1(N1137), .S(N1571), .Z(n428) );
  CMX2X1 U634 ( .A0(\memory[12][2] ), .A1(N1139), .S(N1571), .Z(n427) );
  CMX2X1 U635 ( .A0(\memory[12][3] ), .A1(N1141), .S(N1571), .Z(n426) );
  CMX2X1 U636 ( .A0(\memory[13][0] ), .A1(N1143), .S(N1575), .Z(n425) );
  CMX2X1 U637 ( .A0(\memory[13][1] ), .A1(N1145), .S(N1575), .Z(n424) );
  CMX2X1 U638 ( .A0(\memory[13][2] ), .A1(N1147), .S(N1575), .Z(n423) );
  CMX2X1 U639 ( .A0(\memory[13][3] ), .A1(N1149), .S(N1575), .Z(n422) );
  CMX2X1 U640 ( .A0(\memory[14][0] ), .A1(N1151), .S(N1579), .Z(n421) );
  CMX2X1 U641 ( .A0(\memory[14][1] ), .A1(N1153), .S(N1579), .Z(n420) );
  CMX2X1 U642 ( .A0(\memory[14][2] ), .A1(N1155), .S(N1579), .Z(n419) );
  CMX2X1 U643 ( .A0(\memory[14][3] ), .A1(N1157), .S(N1579), .Z(n418) );
  CMX2X1 U644 ( .A0(\memory[15][0] ), .A1(N1159), .S(N1583), .Z(n417) );
  CMX2X1 U645 ( .A0(\memory[15][1] ), .A1(N1161), .S(N1583), .Z(n416) );
  CMX2X1 U646 ( .A0(\memory[15][2] ), .A1(N1163), .S(N1583), .Z(n415) );
  CMX2X1 U647 ( .A0(\memory[15][3] ), .A1(N1165), .S(N1583), .Z(n414) );
  CMX2X1 U648 ( .A0(\memory[16][0] ), .A1(N1167), .S(N1587), .Z(n413) );
  CMX2X1 U649 ( .A0(\memory[16][1] ), .A1(N1169), .S(N1587), .Z(n412) );
  CMX2X1 U650 ( .A0(\memory[16][2] ), .A1(N1171), .S(N1587), .Z(n411) );
  CMX2X1 U651 ( .A0(\memory[16][3] ), .A1(N1173), .S(N1587), .Z(n410) );
  CMX2X1 U652 ( .A0(\memory[17][0] ), .A1(N1175), .S(N1591), .Z(n409) );
  CMX2X1 U653 ( .A0(\memory[17][1] ), .A1(N1177), .S(N1591), .Z(n408) );
  CMX2X1 U654 ( .A0(\memory[17][2] ), .A1(N1179), .S(N1591), .Z(n407) );
  CMX2X1 U655 ( .A0(\memory[17][3] ), .A1(N1181), .S(N1591), .Z(n406) );
  CMX2X1 U656 ( .A0(\memory[18][0] ), .A1(N1183), .S(N1595), .Z(n405) );
  CMX2X1 U657 ( .A0(\memory[18][1] ), .A1(N1185), .S(N1595), .Z(n404) );
  CMX2X1 U658 ( .A0(\memory[18][2] ), .A1(N1187), .S(N1595), .Z(n403) );
  CMX2X1 U659 ( .A0(\memory[18][3] ), .A1(N1189), .S(N1595), .Z(n402) );
  CMX2X1 U660 ( .A0(\memory[19][0] ), .A1(N1191), .S(N1599), .Z(n401) );
  CMX2X1 U661 ( .A0(\memory[19][1] ), .A1(N1193), .S(N1599), .Z(n400) );
  CMX2X1 U662 ( .A0(\memory[19][2] ), .A1(N1195), .S(N1599), .Z(n399) );
  CMX2X1 U663 ( .A0(\memory[19][3] ), .A1(N1197), .S(N1599), .Z(n398) );
  CMX2X1 U664 ( .A0(\memory[20][0] ), .A1(N1199), .S(N1603), .Z(n397) );
  CMX2X1 U665 ( .A0(\memory[20][1] ), .A1(N1201), .S(N1603), .Z(n396) );
  CMX2X1 U666 ( .A0(\memory[20][2] ), .A1(N1203), .S(N1603), .Z(n395) );
  CMX2X1 U667 ( .A0(\memory[20][3] ), .A1(N1205), .S(N1603), .Z(n394) );
  CMX2X1 U668 ( .A0(\memory[21][0] ), .A1(N1207), .S(N1607), .Z(n393) );
  CMX2X1 U669 ( .A0(\memory[21][1] ), .A1(N1209), .S(N1607), .Z(n392) );
  CMX2X1 U670 ( .A0(\memory[21][2] ), .A1(N1211), .S(N1607), .Z(n391) );
  CMX2X1 U671 ( .A0(\memory[21][3] ), .A1(N1213), .S(N1607), .Z(n390) );
  CMX2X1 U672 ( .A0(\memory[22][0] ), .A1(N1215), .S(N1611), .Z(n389) );
  CMX2X1 U673 ( .A0(\memory[22][1] ), .A1(N1217), .S(N1611), .Z(n388) );
  CMX2X1 U674 ( .A0(\memory[22][2] ), .A1(N1219), .S(N1611), .Z(n387) );
  CMX2X1 U675 ( .A0(\memory[22][3] ), .A1(N1221), .S(N1611), .Z(n386) );
  CMX2X1 U676 ( .A0(\memory[23][0] ), .A1(N1223), .S(N1615), .Z(n385) );
  CMX2X1 U677 ( .A0(\memory[23][1] ), .A1(N1225), .S(N1615), .Z(n384) );
  CMX2X1 U678 ( .A0(\memory[23][2] ), .A1(N1227), .S(N1615), .Z(n383) );
  CMX2X1 U679 ( .A0(\memory[23][3] ), .A1(N1229), .S(N1615), .Z(n382) );
  CMX2X1 U680 ( .A0(\memory[24][0] ), .A1(N1231), .S(N1619), .Z(n381) );
  CMX2X1 U681 ( .A0(\memory[24][1] ), .A1(N1233), .S(N1619), .Z(n380) );
  CMX2X1 U682 ( .A0(\memory[24][2] ), .A1(N1235), .S(N1619), .Z(n379) );
  CMX2X1 U683 ( .A0(\memory[24][3] ), .A1(N1237), .S(N1619), .Z(n378) );
  CMX2X1 U684 ( .A0(\memory[25][0] ), .A1(N1239), .S(N1623), .Z(n377) );
  CMX2X1 U685 ( .A0(\memory[25][1] ), .A1(N1241), .S(N1623), .Z(n376) );
  CMX2X1 U686 ( .A0(\memory[25][2] ), .A1(N1243), .S(N1623), .Z(n375) );
  CMX2X1 U687 ( .A0(\memory[25][3] ), .A1(N1245), .S(N1623), .Z(n374) );
  CMX2X1 U688 ( .A0(\memory[26][0] ), .A1(N1247), .S(N1627), .Z(n373) );
  CMX2X1 U689 ( .A0(\memory[26][1] ), .A1(N1249), .S(N1627), .Z(n372) );
  CMX2X1 U690 ( .A0(\memory[26][2] ), .A1(N1251), .S(N1627), .Z(n371) );
  CMX2X1 U691 ( .A0(\memory[26][3] ), .A1(N1253), .S(N1627), .Z(n370) );
  CMX2X1 U692 ( .A0(\memory[27][0] ), .A1(N1255), .S(N1631), .Z(n369) );
  CMX2X1 U693 ( .A0(\memory[27][1] ), .A1(N1257), .S(N1631), .Z(n368) );
  CMX2X1 U694 ( .A0(\memory[27][2] ), .A1(N1259), .S(N1631), .Z(n367) );
  CMX2X1 U695 ( .A0(\memory[27][3] ), .A1(N1261), .S(N1631), .Z(n366) );
  CMX2X1 U696 ( .A0(\memory[28][0] ), .A1(N1263), .S(N1635), .Z(n365) );
  CMX2X1 U697 ( .A0(\memory[28][1] ), .A1(N1265), .S(N1635), .Z(n364) );
  CMX2X1 U698 ( .A0(\memory[28][2] ), .A1(N1267), .S(N1635), .Z(n363) );
  CMX2X1 U699 ( .A0(\memory[28][3] ), .A1(N1269), .S(N1635), .Z(n362) );
  CMX2X1 U700 ( .A0(\memory[29][0] ), .A1(N1271), .S(N1639), .Z(n361) );
  CMX2X1 U701 ( .A0(\memory[29][1] ), .A1(N1273), .S(N1639), .Z(n360) );
  CMX2X1 U702 ( .A0(\memory[29][2] ), .A1(N1275), .S(N1639), .Z(n359) );
  CMX2X1 U703 ( .A0(\memory[29][3] ), .A1(N1277), .S(N1639), .Z(n358) );
  CMX2X1 U704 ( .A0(\memory[30][0] ), .A1(N1279), .S(N1643), .Z(n357) );
  CMX2X1 U705 ( .A0(\memory[30][1] ), .A1(N1281), .S(N1643), .Z(n356) );
  CMX2X1 U706 ( .A0(\memory[30][2] ), .A1(N1283), .S(N1643), .Z(n355) );
  CMX2X1 U707 ( .A0(\memory[30][3] ), .A1(N1285), .S(N1643), .Z(n354) );
  CMX2X1 U709 ( .A0(full), .A1(n652), .S(N1483), .Z(n352) );
  fifo_DW01_inc_0 add_74 ( .A({N248, N249, N250, N251, N252, N253, N254, N255, 
        N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
        N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279}), .SUM({N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, 
        N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, 
        N571, N570, N569, N568, N567, N566, N565, N564, N563}) );
  fifo_DW01_sub_0 sub_42_aco ( .A({n634, counter[30:27], n614, n613, 
        counter[24:0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        rd_enable}), .CI(1'b0), .DIFF({N123, N121, N119, N117, N115, N113, 
        N111, N109, N107, N105, N103, N101, N99, N97, N95, N93, N91, N89, N87, 
        N85, N83, N81, N79, N77, N75, N73, N71, N69, N67, N65, N63, N61}) );
  CFD2X1 \counter_reg[31]  ( .D(n516), .CP(clock), .CD(reset), .Q(n634), .QN(
        n547) );
  CFD2QX1 \counter_reg[24]  ( .D(n492), .CP(clock), .CD(reset), .Q(counter[24]) );
  CFD2QX1 full_reg ( .D(n352), .CP(clock), .CD(reset), .Q(full) );
  CFD2QX1 \counter_reg[9]  ( .D(n507), .CP(clock), .CD(reset), .Q(counter[9])
         );
  CFD2QX1 \counter_reg[8]  ( .D(n508), .CP(clock), .CD(reset), .Q(counter[8])
         );
  CFD2QX1 \counter_reg[7]  ( .D(n509), .CP(clock), .CD(reset), .Q(counter[7])
         );
  CFD2QX1 \counter_reg[5]  ( .D(n511), .CP(clock), .CD(reset), .Q(counter[5])
         );
  CFD2QX1 \counter_reg[21]  ( .D(n495), .CP(clock), .CD(reset), .Q(counter[21]) );
  CFD2QX1 \counter_reg[20]  ( .D(n496), .CP(clock), .CD(reset), .Q(counter[20]) );
  CFD2QX1 \counter_reg[19]  ( .D(n497), .CP(clock), .CD(reset), .Q(counter[19]) );
  CFD2QX1 \counter_reg[17]  ( .D(n499), .CP(clock), .CD(reset), .Q(counter[17]) );
  CFD2QX1 \counter_reg[14]  ( .D(n502), .CP(clock), .CD(reset), .Q(counter[14]) );
  CFD2QX1 \counter_reg[11]  ( .D(n505), .CP(clock), .CD(reset), .Q(counter[11]) );
  CFD2QX1 \counter_reg[10]  ( .D(n506), .CP(clock), .CD(reset), .Q(counter[10]) );
  CFD2QX1 \counter_reg[6]  ( .D(n510), .CP(clock), .CD(reset), .Q(counter[6])
         );
  CFD2QX1 \counter_reg[18]  ( .D(n498), .CP(clock), .CD(reset), .Q(counter[18]) );
  CFD2QX1 \counter_reg[3]  ( .D(n513), .CP(clock), .CD(reset), .Q(counter[3])
         );
  CFD2QX1 \counter_reg[23]  ( .D(n493), .CP(clock), .CD(reset), .Q(counter[23]) );
  CFD2QX1 \counter_reg[22]  ( .D(n494), .CP(clock), .CD(reset), .Q(counter[22]) );
  CFD2QX1 \counter_reg[12]  ( .D(n504), .CP(clock), .CD(reset), .Q(counter[12]) );
  CFD2QX1 \counter_reg[15]  ( .D(n501), .CP(clock), .CD(reset), .Q(counter[15]) );
  CFD2QX1 \counter_reg[16]  ( .D(n500), .CP(clock), .CD(reset), .Q(counter[16]) );
  CFD2QX1 \counter_reg[13]  ( .D(n503), .CP(clock), .CD(reset), .Q(counter[13]) );
  CFD2QX1 \counter_reg[4]  ( .D(n512), .CP(clock), .CD(reset), .Q(counter[4])
         );
  CFD2QX1 \counter_reg[2]  ( .D(n514), .CP(clock), .CD(reset), .Q(counter[2])
         );
  CFD2QX1 \counter_reg[1]  ( .D(n515), .CP(clock), .CD(reset), .Q(counter[1])
         );
  CFD2QX1 \counter_reg[0]  ( .D(n517), .CP(clock), .CD(reset), .Q(counter[0])
         );
  CFD2QX1 \counter_reg[25]  ( .D(n491), .CP(clock), .CD(reset), .Q(n607) );
  CFD2QX1 \counter_reg[26]  ( .D(n490), .CP(clock), .CD(reset), .Q(n609) );
  CFD2QX1 \counter_reg[27]  ( .D(n489), .CP(clock), .CD(reset), .Q(counter[27]) );
  CFD2QX1 \counter_reg[28]  ( .D(n488), .CP(clock), .CD(reset), .Q(counter[28]) );
  CFD2QX1 \counter_reg[30]  ( .D(n486), .CP(clock), .CD(reset), .Q(counter[30]) );
  CFD2QX1 \counter_reg[29]  ( .D(n487), .CP(clock), .CD(reset), .Q(counter[29]) );
  CFD1QXL \code_reg[3]  ( .D(n474), .CP(clock), .Q(code[3]) );
  CFD1QXL \code_reg[2]  ( .D(n476), .CP(clock), .Q(code[2]) );
  CFD1QXL \code_reg[1]  ( .D(n478), .CP(clock), .Q(code[1]) );
  CFD1QXL \code_reg[0]  ( .D(n480), .CP(clock), .Q(code[0]) );
  CFD1QXL \memory_reg[31][3]  ( .D(n520), .CP(clock), .Q(\memory[31][3] ) );
  CFD1QXL \memory_reg[31][2]  ( .D(n523), .CP(clock), .Q(\memory[31][2] ) );
  CFD1QXL \memory_reg[31][1]  ( .D(n526), .CP(clock), .Q(\memory[31][1] ) );
  CFD1QXL \memory_reg[31][0]  ( .D(n529), .CP(clock), .Q(\memory[31][0] ) );
  CFD1QXL \memory_reg[30][2]  ( .D(n355), .CP(clock), .Q(\memory[30][2] ) );
  CFD1QXL \memory_reg[30][0]  ( .D(n357), .CP(clock), .Q(\memory[30][0] ) );
  CFD1QXL \memory_reg[29][2]  ( .D(n359), .CP(clock), .Q(\memory[29][2] ) );
  CFD1QXL \memory_reg[29][0]  ( .D(n361), .CP(clock), .Q(\memory[29][0] ) );
  CFD1QXL \memory_reg[28][2]  ( .D(n363), .CP(clock), .Q(\memory[28][2] ) );
  CFD1QXL \memory_reg[28][0]  ( .D(n365), .CP(clock), .Q(\memory[28][0] ) );
  CFD1QXL \memory_reg[27][2]  ( .D(n367), .CP(clock), .Q(\memory[27][2] ) );
  CFD1QXL \memory_reg[27][0]  ( .D(n369), .CP(clock), .Q(\memory[27][0] ) );
  CFD1QXL \memory_reg[26][2]  ( .D(n371), .CP(clock), .Q(\memory[26][2] ) );
  CFD1QXL \memory_reg[26][0]  ( .D(n373), .CP(clock), .Q(\memory[26][0] ) );
  CFD1QXL \memory_reg[25][2]  ( .D(n375), .CP(clock), .Q(\memory[25][2] ) );
  CFD1QXL \memory_reg[25][0]  ( .D(n377), .CP(clock), .Q(\memory[25][0] ) );
  CFD1QXL \memory_reg[24][2]  ( .D(n379), .CP(clock), .Q(\memory[24][2] ) );
  CFD1QXL \memory_reg[24][0]  ( .D(n381), .CP(clock), .Q(\memory[24][0] ) );
  CFD1QXL \memory_reg[23][2]  ( .D(n383), .CP(clock), .Q(\memory[23][2] ) );
  CFD1QXL \memory_reg[23][0]  ( .D(n385), .CP(clock), .Q(\memory[23][0] ) );
  CFD1QXL \memory_reg[22][2]  ( .D(n387), .CP(clock), .Q(\memory[22][2] ) );
  CFD1QXL \memory_reg[22][0]  ( .D(n389), .CP(clock), .Q(\memory[22][0] ) );
  CFD1QXL \memory_reg[21][2]  ( .D(n391), .CP(clock), .Q(\memory[21][2] ) );
  CFD1QXL \memory_reg[21][0]  ( .D(n393), .CP(clock), .Q(\memory[21][0] ) );
  CFD1QXL \memory_reg[20][2]  ( .D(n395), .CP(clock), .Q(\memory[20][2] ) );
  CFD1QXL \memory_reg[20][0]  ( .D(n397), .CP(clock), .Q(\memory[20][0] ) );
  CFD1QXL \memory_reg[19][2]  ( .D(n399), .CP(clock), .Q(\memory[19][2] ) );
  CFD1QXL \memory_reg[19][0]  ( .D(n401), .CP(clock), .Q(\memory[19][0] ) );
  CFD1QXL \memory_reg[18][2]  ( .D(n403), .CP(clock), .Q(\memory[18][2] ) );
  CFD1QXL \memory_reg[18][0]  ( .D(n405), .CP(clock), .Q(\memory[18][0] ) );
  CFD1QXL \memory_reg[17][2]  ( .D(n407), .CP(clock), .Q(\memory[17][2] ) );
  CFD1QXL \memory_reg[17][0]  ( .D(n409), .CP(clock), .Q(\memory[17][0] ) );
  CFD1QXL \memory_reg[16][2]  ( .D(n411), .CP(clock), .Q(\memory[16][2] ) );
  CFD1QXL \memory_reg[16][0]  ( .D(n413), .CP(clock), .Q(\memory[16][0] ) );
  CFD1QXL \memory_reg[15][2]  ( .D(n415), .CP(clock), .Q(\memory[15][2] ) );
  CFD1QXL \memory_reg[15][0]  ( .D(n417), .CP(clock), .Q(\memory[15][0] ) );
  CFD1QXL \memory_reg[14][2]  ( .D(n419), .CP(clock), .Q(\memory[14][2] ) );
  CFD1QXL \memory_reg[14][0]  ( .D(n421), .CP(clock), .Q(\memory[14][0] ) );
  CFD1QXL \memory_reg[13][2]  ( .D(n423), .CP(clock), .Q(\memory[13][2] ) );
  CFD1QXL \memory_reg[13][0]  ( .D(n425), .CP(clock), .Q(\memory[13][0] ) );
  CFD1QXL \memory_reg[12][2]  ( .D(n427), .CP(clock), .Q(\memory[12][2] ) );
  CFD1QXL \memory_reg[12][0]  ( .D(n429), .CP(clock), .Q(\memory[12][0] ) );
  CFD1QXL \memory_reg[11][2]  ( .D(n431), .CP(clock), .Q(\memory[11][2] ) );
  CFD1QXL \memory_reg[11][0]  ( .D(n433), .CP(clock), .Q(\memory[11][0] ) );
  CFD1QXL \memory_reg[10][2]  ( .D(n435), .CP(clock), .Q(\memory[10][2] ) );
  CFD1QXL \memory_reg[10][0]  ( .D(n437), .CP(clock), .Q(\memory[10][0] ) );
  CFD1QXL \memory_reg[9][2]  ( .D(n439), .CP(clock), .Q(\memory[9][2] ) );
  CFD1QXL \memory_reg[9][0]  ( .D(n441), .CP(clock), .Q(\memory[9][0] ) );
  CFD1QXL \memory_reg[8][2]  ( .D(n443), .CP(clock), .Q(\memory[8][2] ) );
  CFD1QXL \memory_reg[8][0]  ( .D(n445), .CP(clock), .Q(\memory[8][0] ) );
  CFD1QXL \memory_reg[7][2]  ( .D(n447), .CP(clock), .Q(\memory[7][2] ) );
  CFD1QXL \memory_reg[7][0]  ( .D(n449), .CP(clock), .Q(\memory[7][0] ) );
  CFD1QXL \memory_reg[6][2]  ( .D(n451), .CP(clock), .Q(\memory[6][2] ) );
  CFD1QXL \memory_reg[6][0]  ( .D(n453), .CP(clock), .Q(\memory[6][0] ) );
  CFD1QXL \memory_reg[5][2]  ( .D(n455), .CP(clock), .Q(\memory[5][2] ) );
  CFD1QXL \memory_reg[5][0]  ( .D(n457), .CP(clock), .Q(\memory[5][0] ) );
  CFD1QXL \memory_reg[4][2]  ( .D(n459), .CP(clock), .Q(\memory[4][2] ) );
  CFD1QXL \memory_reg[4][0]  ( .D(n461), .CP(clock), .Q(\memory[4][0] ) );
  CFD1QXL \memory_reg[3][2]  ( .D(n463), .CP(clock), .Q(\memory[3][2] ) );
  CFD1QXL \memory_reg[3][0]  ( .D(n465), .CP(clock), .Q(\memory[3][0] ) );
  CFD1QXL \memory_reg[2][2]  ( .D(n467), .CP(clock), .Q(\memory[2][2] ) );
  CFD1QXL \memory_reg[2][0]  ( .D(n469), .CP(clock), .Q(\memory[2][0] ) );
  CFD1QXL \memory_reg[1][2]  ( .D(n471), .CP(clock), .Q(\memory[1][2] ) );
  CFD1QXL \memory_reg[1][0]  ( .D(n473), .CP(clock), .Q(\memory[1][0] ) );
  CFD1QXL \memory_reg[0][2]  ( .D(n477), .CP(clock), .Q(\memory[0][2] ) );
  CFD1QXL \memory_reg[0][0]  ( .D(n481), .CP(clock), .Q(\memory[0][0] ) );
  CFD1QXL \memory_reg[29][3]  ( .D(n358), .CP(clock), .Q(\memory[29][3] ) );
  CFD1QXL \memory_reg[29][1]  ( .D(n360), .CP(clock), .Q(\memory[29][1] ) );
  CFD1QXL \memory_reg[28][3]  ( .D(n362), .CP(clock), .Q(\memory[28][3] ) );
  CFD1QXL \memory_reg[28][1]  ( .D(n364), .CP(clock), .Q(\memory[28][1] ) );
  CFD1QXL \memory_reg[27][3]  ( .D(n366), .CP(clock), .Q(\memory[27][3] ) );
  CFD1QXL \memory_reg[27][1]  ( .D(n368), .CP(clock), .Q(\memory[27][1] ) );
  CFD1QXL \memory_reg[26][3]  ( .D(n370), .CP(clock), .Q(\memory[26][3] ) );
  CFD1QXL \memory_reg[26][1]  ( .D(n372), .CP(clock), .Q(\memory[26][1] ) );
  CFD1QXL \memory_reg[25][3]  ( .D(n374), .CP(clock), .Q(\memory[25][3] ) );
  CFD1QXL \memory_reg[25][1]  ( .D(n376), .CP(clock), .Q(\memory[25][1] ) );
  CFD1QXL \memory_reg[24][3]  ( .D(n378), .CP(clock), .Q(\memory[24][3] ) );
  CFD1QXL \memory_reg[24][1]  ( .D(n380), .CP(clock), .Q(\memory[24][1] ) );
  CFD1QXL \memory_reg[23][3]  ( .D(n382), .CP(clock), .Q(\memory[23][3] ) );
  CFD1QXL \memory_reg[23][1]  ( .D(n384), .CP(clock), .Q(\memory[23][1] ) );
  CFD1QXL \memory_reg[22][3]  ( .D(n386), .CP(clock), .Q(\memory[22][3] ) );
  CFD1QXL \memory_reg[22][1]  ( .D(n388), .CP(clock), .Q(\memory[22][1] ) );
  CFD1QXL \memory_reg[21][3]  ( .D(n390), .CP(clock), .Q(\memory[21][3] ) );
  CFD1QXL \memory_reg[21][1]  ( .D(n392), .CP(clock), .Q(\memory[21][1] ) );
  CFD1QXL \memory_reg[20][3]  ( .D(n394), .CP(clock), .Q(\memory[20][3] ) );
  CFD1QXL \memory_reg[20][1]  ( .D(n396), .CP(clock), .Q(\memory[20][1] ) );
  CFD1QXL \memory_reg[19][3]  ( .D(n398), .CP(clock), .Q(\memory[19][3] ) );
  CFD1QXL \memory_reg[19][1]  ( .D(n400), .CP(clock), .Q(\memory[19][1] ) );
  CFD1QXL \memory_reg[18][3]  ( .D(n402), .CP(clock), .Q(\memory[18][3] ) );
  CFD1QXL \memory_reg[18][1]  ( .D(n404), .CP(clock), .Q(\memory[18][1] ) );
  CFD1QXL \memory_reg[17][3]  ( .D(n406), .CP(clock), .Q(\memory[17][3] ) );
  CFD1QXL \memory_reg[17][1]  ( .D(n408), .CP(clock), .Q(\memory[17][1] ) );
  CFD1QXL \memory_reg[16][3]  ( .D(n410), .CP(clock), .Q(\memory[16][3] ) );
  CFD1QXL \memory_reg[16][1]  ( .D(n412), .CP(clock), .Q(\memory[16][1] ) );
  CFD1QXL \memory_reg[15][3]  ( .D(n414), .CP(clock), .Q(\memory[15][3] ) );
  CFD1QXL \memory_reg[15][1]  ( .D(n416), .CP(clock), .Q(\memory[15][1] ) );
  CFD1QXL \memory_reg[14][3]  ( .D(n418), .CP(clock), .Q(\memory[14][3] ) );
  CFD1QXL \memory_reg[14][1]  ( .D(n420), .CP(clock), .Q(\memory[14][1] ) );
  CFD1QXL \memory_reg[13][3]  ( .D(n422), .CP(clock), .Q(\memory[13][3] ) );
  CFD1QXL \memory_reg[13][1]  ( .D(n424), .CP(clock), .Q(\memory[13][1] ) );
  CFD1QXL \memory_reg[12][3]  ( .D(n426), .CP(clock), .Q(\memory[12][3] ) );
  CFD1QXL \memory_reg[12][1]  ( .D(n428), .CP(clock), .Q(\memory[12][1] ) );
  CFD1QXL \memory_reg[11][3]  ( .D(n430), .CP(clock), .Q(\memory[11][3] ) );
  CFD1QXL \memory_reg[11][1]  ( .D(n432), .CP(clock), .Q(\memory[11][1] ) );
  CFD1QXL \memory_reg[10][3]  ( .D(n434), .CP(clock), .Q(\memory[10][3] ) );
  CFD1QXL \memory_reg[10][1]  ( .D(n436), .CP(clock), .Q(\memory[10][1] ) );
  CFD1QXL \memory_reg[9][3]  ( .D(n438), .CP(clock), .Q(\memory[9][3] ) );
  CFD1QXL \memory_reg[9][1]  ( .D(n440), .CP(clock), .Q(\memory[9][1] ) );
  CFD1QXL \memory_reg[8][3]  ( .D(n442), .CP(clock), .Q(\memory[8][3] ) );
  CFD1QXL \memory_reg[8][1]  ( .D(n444), .CP(clock), .Q(\memory[8][1] ) );
  CFD1QXL \memory_reg[7][3]  ( .D(n446), .CP(clock), .Q(\memory[7][3] ) );
  CFD1QXL \memory_reg[7][1]  ( .D(n448), .CP(clock), .Q(\memory[7][1] ) );
  CFD1QXL \memory_reg[6][3]  ( .D(n450), .CP(clock), .Q(\memory[6][3] ) );
  CFD1QXL \memory_reg[6][1]  ( .D(n452), .CP(clock), .Q(\memory[6][1] ) );
  CFD1QXL \memory_reg[5][3]  ( .D(n454), .CP(clock), .Q(\memory[5][3] ) );
  CFD1QXL \memory_reg[5][1]  ( .D(n456), .CP(clock), .Q(\memory[5][1] ) );
  CFD1QXL \memory_reg[4][3]  ( .D(n458), .CP(clock), .Q(\memory[4][3] ) );
  CFD1QXL \memory_reg[4][1]  ( .D(n460), .CP(clock), .Q(\memory[4][1] ) );
  CFD1QXL \memory_reg[3][3]  ( .D(n462), .CP(clock), .Q(\memory[3][3] ) );
  CFD1QXL \memory_reg[3][1]  ( .D(n464), .CP(clock), .Q(\memory[3][1] ) );
  CFD1QXL \memory_reg[2][3]  ( .D(n466), .CP(clock), .Q(\memory[2][3] ) );
  CFD1QXL \memory_reg[2][1]  ( .D(n468), .CP(clock), .Q(\memory[2][1] ) );
  CFD1QXL \memory_reg[1][3]  ( .D(n470), .CP(clock), .Q(\memory[1][3] ) );
  CFD1QXL \memory_reg[1][1]  ( .D(n472), .CP(clock), .Q(\memory[1][1] ) );
  CFD1QXL \memory_reg[0][3]  ( .D(n475), .CP(clock), .Q(\memory[0][3] ) );
  CIVXL U710 ( .A(reset), .Z(n14) );
  CNIVXL U711 ( .A(wr_enable), .Z(n518) );
  CNIVX1 U712 ( .A(\memory[0][1] ), .Z(n519) );
  CAN2XL U713 ( .A(n657), .B(reset), .Z(N1651) );
  CMX2X4 U714 ( .A0(\memory[31][3] ), .A1(data[3]), .S(N1647), .Z(n482) );
  CNIVX1 U715 ( .A(n521), .Z(n520) );
  CNIVX1 U716 ( .A(n522), .Z(n521) );
  CNIVX1 U717 ( .A(n482), .Z(n522) );
  CMX2X4 U718 ( .A0(\memory[31][2] ), .A1(data[2]), .S(N1647), .Z(n483) );
  CNIVX1 U719 ( .A(n524), .Z(n523) );
  CNIVX1 U720 ( .A(n525), .Z(n524) );
  CNIVX1 U721 ( .A(n483), .Z(n525) );
  CMX2X4 U722 ( .A0(\memory[31][1] ), .A1(data[1]), .S(N1647), .Z(n484) );
  CNIVX1 U723 ( .A(n527), .Z(n526) );
  CNIVX1 U724 ( .A(n528), .Z(n527) );
  CNIVX1 U725 ( .A(n484), .Z(n528) );
  CMX2X4 U726 ( .A0(\memory[31][0] ), .A1(data[0]), .S(N1647), .Z(n485) );
  CNIVX1 U727 ( .A(n530), .Z(n529) );
  CNIVX1 U728 ( .A(n531), .Z(n530) );
  CNIVX1 U729 ( .A(n485), .Z(n531) );
  CANR2XL U730 ( .A(N113), .B(n652), .C(N589), .D(n18), .Z(n27) );
  CAOR2XL U731 ( .A(n76), .B(N1702), .C(\memory[31][3] ), .D(n77), .Z(N1285)
         );
  CAN2X1 U732 ( .A(n589), .B(N113), .Z(N1748) );
  CANR2XL U733 ( .A(N117), .B(n652), .C(N591), .D(n18), .Z(n23) );
  CAOR2XL U734 ( .A(n79), .B(N1702), .C(\memory[31][1] ), .D(n77), .Z(N1281)
         );
  CAN2X1 U735 ( .A(n572), .B(N117), .Z(N1742) );
  CIVXL U736 ( .A(n559), .Z(n564) );
  CIVDX1 U737 ( .A(n557), .Z0(n581), .Z1(n582) );
  COR2X1 U738 ( .A(n533), .B(N1037), .Z(n532) );
  CIVX20 U739 ( .A(n532), .Z(n80) );
  CIVX20 U740 ( .A(data[0]), .Z(n533) );
  COND4CXL U741 ( .A(n605), .B(n681), .C(n680), .D(n679), .Z(n683) );
  CMX2XL U742 ( .A0(counter[0]), .A1(N1291), .S(N1519), .Z(n517) );
  CNR2X1 U743 ( .A(N1682), .B(counter[0]), .Z(n639) );
  CNR5XL U744 ( .A(counter[0]), .B(n678), .C(counter[1]), .D(counter[3]), .E(
        counter[2]), .Z(n680) );
  CNR2IX2 U745 ( .B(data[2]), .A(N1037), .Z(n78) );
  CND2X2 U746 ( .A(N282), .B(n518), .Z(N1037) );
  CND2X1 U747 ( .A(n575), .B(counter[3]), .Z(n554) );
  CDLY1X2 U748 ( .A(N1035), .Z(n641) );
  CDLY1X2 U749 ( .A(N1035), .Z(n642) );
  CDLY1X2 U750 ( .A(N1035), .Z(n643) );
  CDLY1X2 U751 ( .A(N1035), .Z(n644) );
  CDLY1X2 U752 ( .A(N1035), .Z(n645) );
  CDLY1X2 U753 ( .A(N1035), .Z(n646) );
  CDLY1X2 U754 ( .A(N1035), .Z(n647) );
  CDLY1X2 U755 ( .A(N1035), .Z(n648) );
  CDLY1X2 U756 ( .A(N1035), .Z(n649) );
  CDLY1X2 U757 ( .A(N1035), .Z(n651) );
  CDLY1X2 U758 ( .A(N1035), .Z(n650) );
  CAN2X1 U759 ( .A(n568), .B(N121), .Z(N1736) );
  CMX2XL U760 ( .A0(empty), .A1(N1037), .S(N1482), .Z(n353) );
  CND2X2 U761 ( .A(n551), .B(n550), .Z(N279) );
  CAN2XL U762 ( .A(N276), .B(N1), .Z(N1686) );
  CAN2XL U763 ( .A(N276), .B(N275), .Z(N1684) );
  CAN2XL U764 ( .A(n575), .B(counter[21]), .Z(N1765) );
  CIVX1 U765 ( .A(n560), .Z(n575) );
  CAN2XL U766 ( .A(n552), .B(N3), .Z(N1687) );
  CAN2XL U767 ( .A(n552), .B(N275), .Z(N1685) );
  CIVX1 U768 ( .A(n610), .Z(n614) );
  CMX2X1 U769 ( .A0(n614), .A1(N1343), .S(N1519), .Z(n490) );
  CIVX1 U770 ( .A(n558), .Z(n574) );
  CIVDX2 U771 ( .A(n15), .Z0(n558), .Z1(n559) );
  CND2XL U772 ( .A(N252), .B(n13), .Z(n26) );
  CANR2XL U773 ( .A(N115), .B(n652), .C(N590), .D(n18), .Z(n25) );
  CAN2X1 U774 ( .A(n571), .B(N115), .Z(N1745) );
  CND2IX1 U775 ( .B(n534), .A(n541), .Z(n486) );
  CAN2XL U776 ( .A(counter[30]), .B(n540), .Z(n534) );
  CND2X1 U777 ( .A(N593), .B(n18), .Z(n546) );
  CND2X1 U778 ( .A(N1351), .B(N1519), .Z(n541) );
  CND2X2 U779 ( .A(N594), .B(n18), .Z(n535) );
  COR6X1 U780 ( .A(counter[29]), .B(counter[28]), .C(counter[27]), .D(
        counter[9]), .E(counter[8]), .F(counter[30]), .Z(n686) );
  CND2XL U781 ( .A(N250), .B(n13), .Z(n22) );
  CAN2X1 U782 ( .A(n535), .B(n536), .Z(n548) );
  CAN2X1 U783 ( .A(n537), .B(n542), .Z(n536) );
  CIVX2 U784 ( .A(n544), .Z(n537) );
  CNR2IX1 U785 ( .B(n547), .A(n539), .Z(n538) );
  CNR8X1 U786 ( .A(n685), .B(counter[22]), .C(counter[21]), .D(n614), .E(n613), 
        .F(counter[24]), .G(n686), .H(counter[23]), .Z(n539) );
  CIVXL U787 ( .A(N1519), .Z(n540) );
  CND2XL U788 ( .A(N123), .B(n652), .Z(n542) );
  CNIVX2 U789 ( .A(N1035), .Z(n652) );
  CIVX1 U790 ( .A(n608), .Z(n613) );
  CIVX2 U791 ( .A(n547), .Z(n543) );
  CAN2XL U792 ( .A(n598), .B(counter[23]), .Z(N1759) );
  CAN2XL U793 ( .A(N248), .B(n13), .Z(n544) );
  CIVX2 U794 ( .A(n607), .Z(n608) );
  CMX2XL U795 ( .A0(counter[24]), .A1(N1339), .S(N1519), .Z(n492) );
  CAN2XL U796 ( .A(n597), .B(counter[24]), .Z(N1756) );
  CMX2XL U797 ( .A0(counter[23]), .A1(N1337), .S(N1519), .Z(n493) );
  CND2XL U798 ( .A(N121), .B(n652), .Z(n545) );
  CAN2X1 U799 ( .A(n545), .B(n546), .Z(n19) );
  CAN2XL U800 ( .A(n577), .B(counter[29]), .Z(N1741) );
  CMXI2X1 U801 ( .A0(n547), .A1(n548), .S(N1519), .Z(n516) );
  CND2X1 U802 ( .A(n564), .B(N61), .Z(n550) );
  CIVDXL U803 ( .A(N277), .Z0(N1688) );
  CMX2XL U804 ( .A0(counter[6]), .A1(N1303), .S(N1519), .Z(n510) );
  CAN2XL U805 ( .A(n578), .B(counter[6]), .Z(N1810) );
  CND2X1 U806 ( .A(n573), .B(counter[1]), .Z(n556) );
  CAN2XL U807 ( .A(n573), .B(counter[18]), .Z(N1774) );
  CIVX2 U808 ( .A(n558), .Z(n573) );
  CND2XL U809 ( .A(n15), .B(counter[0]), .Z(n551) );
  CANR2XL U810 ( .A(N85), .B(n651), .C(N575), .D(n18), .Z(n55) );
  CANR2XL U811 ( .A(N87), .B(n651), .C(N576), .D(n18), .Z(n53) );
  CND2XL U812 ( .A(n55), .B(n56), .Z(N1315) );
  CANR2XL U813 ( .A(N91), .B(n651), .C(N578), .D(n18), .Z(n49) );
  CANR2XL U814 ( .A(N93), .B(n651), .C(N579), .D(n18), .Z(n47) );
  CND2XL U815 ( .A(n49), .B(n50), .Z(N1321) );
  CIVXL U816 ( .A(N279), .Z(N4) );
  CIVXL U817 ( .A(N279), .Z(N6) );
  CND2IX2 U818 ( .B(N1823), .A(n556), .Z(N278) );
  CAN2X2 U819 ( .A(n553), .B(n554), .Z(n552) );
  CIVX4 U820 ( .A(n552), .Z(N276) );
  CND2XL U821 ( .A(n567), .B(N67), .Z(n553) );
  CAN2X1 U822 ( .A(N6), .B(N7), .Z(N1692) );
  CANR2XL U823 ( .A(N63), .B(n650), .C(N564), .D(n18), .Z(n74) );
  CANR2XL U824 ( .A(N61), .B(n650), .C(N563), .D(n18), .Z(n75) );
  CANR2XL U825 ( .A(N65), .B(n650), .C(N565), .D(n18), .Z(n73) );
  CND2IX2 U826 ( .B(counter[30]), .A(n632), .Z(N1654) );
  CND2IX2 U827 ( .B(counter[5]), .A(n637), .Z(N1678) );
  CAN2XL U828 ( .A(N279), .B(N7), .Z(N1691) );
  CIVX1 U829 ( .A(n682), .Z(n678) );
  CND2IX1 U830 ( .B(N1820), .A(n555), .Z(N277) );
  CND2XL U831 ( .A(n574), .B(counter[2]), .Z(n555) );
  CANR2XL U832 ( .A(N69), .B(n650), .C(N567), .D(n18), .Z(n71) );
  CAN2XL U833 ( .A(N277), .B(N1692), .Z(N1696) );
  CAN2XL U834 ( .A(N277), .B(N1691), .Z(N1695) );
  CAN2XL U835 ( .A(N277), .B(N1690), .Z(N1694) );
  CAN2XL U836 ( .A(N277), .B(N1689), .Z(N1693) );
  CIVXL U837 ( .A(N278), .Z(N7) );
  CIVX4 U838 ( .A(N98), .Z(n557) );
  CIVDXL U839 ( .A(n15), .Z0(n560), .Z1(n561) );
  CIVDXL U840 ( .A(n15), .Z0(n562), .Z1(n563) );
  CIVX1 U841 ( .A(n559), .Z(n565) );
  CIVX1 U842 ( .A(n559), .Z(n566) );
  CIVXL U843 ( .A(n561), .Z(n567) );
  CIVXL U844 ( .A(n561), .Z(n568) );
  CIVXL U845 ( .A(n561), .Z(n569) );
  CIVXL U846 ( .A(n563), .Z(n570) );
  CIVXL U847 ( .A(n563), .Z(n571) );
  CIVXL U848 ( .A(n563), .Z(n572) );
  CIVXL U849 ( .A(n560), .Z(n576) );
  CIVXL U850 ( .A(n560), .Z(n577) );
  CIVXL U851 ( .A(n562), .Z(n578) );
  CIVXL U852 ( .A(n562), .Z(n579) );
  CIVXL U853 ( .A(n562), .Z(n580) );
  CIVDX1 U854 ( .A(n557), .Z0(n583), .Z1(n584) );
  CIVDXL U855 ( .A(n557), .Z0(n585), .Z1(n586) );
  CIVX1 U856 ( .A(n582), .Z(n587) );
  CIVX1 U857 ( .A(n582), .Z(n588) );
  CIVX1 U858 ( .A(n582), .Z(n589) );
  CIVX2 U859 ( .A(n584), .Z(n590) );
  CIVX2 U860 ( .A(n584), .Z(n591) );
  CIVX2 U861 ( .A(n584), .Z(n592) );
  CIVX2 U862 ( .A(n586), .Z(n593) );
  CIVX2 U863 ( .A(n586), .Z(n594) );
  CIVX2 U864 ( .A(n586), .Z(n595) );
  CIVX1 U865 ( .A(n581), .Z(n596) );
  CIVX1 U866 ( .A(n581), .Z(n597) );
  CIVX1 U867 ( .A(n581), .Z(n598) );
  CIVX2 U868 ( .A(n583), .Z(n599) );
  CIVX2 U869 ( .A(n583), .Z(n600) );
  CIVX2 U870 ( .A(n583), .Z(n601) );
  CIVX2 U871 ( .A(n585), .Z(n602) );
  CIVX2 U872 ( .A(n585), .Z(n603) );
  CIVX2 U873 ( .A(n585), .Z(n604) );
  CIVXL U874 ( .A(n15), .Z(N98) );
  CANR3XL U875 ( .A(counter[5]), .B(counter[4]), .C(counter[7]), .D(counter[6]), .Z(n605) );
  CANR3X2 U876 ( .A(counter[5]), .B(counter[4]), .C(counter[7]), .D(counter[6]), .Z(n682) );
  CND2IX1 U877 ( .B(n609), .A(n608), .Z(n629) );
  CDLY1XL U878 ( .A(n609), .Z(n606) );
  CIVX1 U879 ( .A(n625), .Z(n626) );
  CIVXL U880 ( .A(n606), .Z(n610) );
  CIVX2 U881 ( .A(n623), .Z(n611) );
  CND2IX1 U882 ( .B(N1656), .A(n612), .Z(n620) );
  CNR2X2 U883 ( .A(n615), .B(n611), .Z(n612) );
  CMX2XL U884 ( .A0(counter[22]), .A1(N1335), .S(N1519), .Z(n494) );
  CIVX2 U885 ( .A(counter[22]), .Z(n624) );
  CAN2XL U886 ( .A(n574), .B(counter[22]), .Z(N1762) );
  CMX2XL U887 ( .A0(n613), .A1(N1341), .S(N1519), .Z(n491) );
  CAN2XL U888 ( .A(n579), .B(n613), .Z(N1753) );
  CMX2XL U889 ( .A0(counter[18]), .A1(N1327), .S(N1519), .Z(n498) );
  CAN2X1 U890 ( .A(n599), .B(n614), .Z(N1750) );
  CND2IX1 U891 ( .B(n616), .A(n624), .Z(n615) );
  CND2IX1 U892 ( .B(n629), .A(n622), .Z(n616) );
  CIVX2 U893 ( .A(n619), .Z(n617) );
  CND2IX1 U894 ( .B(n620), .A(n618), .Z(N1667) );
  CNR2X1 U895 ( .A(n621), .B(n617), .Z(n618) );
  CNR2X2 U896 ( .A(counter[17]), .B(counter[16]), .Z(n619) );
  COR2XL U897 ( .A(counter[18]), .B(counter[21]), .Z(n621) );
  CNR2X2 U898 ( .A(counter[24]), .B(counter[23]), .Z(n622) );
  CNR2X2 U899 ( .A(counter[20]), .B(counter[19]), .Z(n623) );
  COR2XL U900 ( .A(counter[10]), .B(counter[9]), .Z(n625) );
  CND2IX1 U901 ( .B(N1672), .A(n626), .Z(N1674) );
  COR2XL U902 ( .A(counter[2]), .B(counter[1]), .Z(n627) );
  CND2IX1 U903 ( .B(N1680), .A(n628), .Z(N1682) );
  CIVX20 U904 ( .A(n627), .Z(n628) );
  CNR2X2 U905 ( .A(counter[28]), .B(N1654), .Z(n630) );
  CND2IX2 U906 ( .B(counter[7]), .A(n636), .Z(n631) );
  CND2IX1 U907 ( .B(counter[27]), .A(n630), .Z(N1656) );
  CNR2X2 U908 ( .A(n631), .B(counter[6]), .Z(n637) );
  CMX2XL U909 ( .A0(counter[29]), .A1(N1349), .S(N1519), .Z(n487) );
  CND2IX2 U910 ( .B(counter[14]), .A(n640), .Z(N1669) );
  CND2IX1 U911 ( .B(counter[11]), .A(n635), .Z(N1672) );
  CNR2X2 U912 ( .A(n634), .B(counter[29]), .Z(n632) );
  COR2XL U913 ( .A(counter[13]), .B(counter[12]), .Z(n633) );
  CNR2X2 U914 ( .A(N1669), .B(n633), .Z(n635) );
  CNR2X2 U915 ( .A(N1674), .B(counter[8]), .Z(n636) );
  CNR2X2 U916 ( .A(N1678), .B(counter[4]), .Z(n638) );
  CND2IX1 U917 ( .B(counter[3]), .A(n638), .Z(N1680) );
  CAN2XL U918 ( .A(n576), .B(counter[30]), .Z(N1738) );
  CNR2X2 U919 ( .A(n639), .B(n538), .Z(N51) );
  CNR2X2 U920 ( .A(N1667), .B(counter[15]), .Z(n640) );
  CAN2XL U921 ( .A(n600), .B(n543), .Z(N1735) );
  CAN2XL U922 ( .A(N4), .B(N278), .Z(N1690) );
  CAN2XL U923 ( .A(N279), .B(N278), .Z(N1689) );
  CAN2XL U924 ( .A(N51), .B(rd_enable), .Z(N247) );
  CNR2IX4 U925 ( .B(rd_enable), .A(N51), .Z(n15) );
  CANR1X4 U926 ( .A(n601), .B(n652), .C(n14), .Z(N1519) );
  CIVXL U927 ( .A(n672), .Z(n653) );
  CIVXL U928 ( .A(n672), .Z(n654) );
  CIVXL U929 ( .A(n672), .Z(n655) );
  CIVXL U930 ( .A(n672), .Z(n656) );
  CIVXL U931 ( .A(n672), .Z(n657) );
  CIVXL U932 ( .A(n672), .Z(n658) );
  CIVXL U933 ( .A(n672), .Z(n659) );
  CIVXL U934 ( .A(n672), .Z(n660) );
  CIVXL U935 ( .A(n672), .Z(n661) );
  CIVXL U936 ( .A(n672), .Z(n662) );
  CNIVX3 U937 ( .A(n677), .Z(n663) );
  CNIVX3 U938 ( .A(n677), .Z(n664) );
  CNIVX3 U939 ( .A(n676), .Z(n665) );
  CNIVX3 U940 ( .A(n676), .Z(n666) );
  CNIVX3 U941 ( .A(n675), .Z(n667) );
  CNIVX3 U942 ( .A(n675), .Z(n668) );
  CNIVX3 U943 ( .A(n674), .Z(n669) );
  CNIVX3 U944 ( .A(n674), .Z(n670) );
  CNIVX3 U945 ( .A(n673), .Z(n671) );
  CNIVX3 U946 ( .A(n673), .Z(n672) );
  CIVX2 U947 ( .A(N247), .Z(n673) );
  CIVX2 U948 ( .A(N247), .Z(n674) );
  CIVX2 U949 ( .A(N247), .Z(n675) );
  CIVX2 U950 ( .A(N247), .Z(n676) );
  CIVX2 U951 ( .A(N247), .Z(n677) );
  COR3X1 U952 ( .A(counter[14]), .B(counter[13]), .C(counter[12]), .Z(n684) );
  CIVX1 U953 ( .A(counter[5]), .Z(n681) );
  CNR2X1 U954 ( .A(counter[11]), .B(counter[10]), .Z(n679) );
  COR8X1 U955 ( .A(counter[17]), .B(counter[16]), .C(counter[15]), .D(
        counter[20]), .E(counter[19]), .F(counter[18]), .G(n684), .H(n683), 
        .Z(n685) );
  COR6X1 U956 ( .A(N267), .B(N268), .C(N269), .D(N264), .E(N265), .F(N266), 
        .Z(n687) );
  CNR8X1 U957 ( .A(n687), .B(N263), .C(N261), .D(N262), .E(N257), .F(N258), 
        .G(N259), .H(N260), .Z(n690) );
  COR6X1 U958 ( .A(N254), .B(N255), .C(N256), .D(N251), .E(N252), .F(N253), 
        .Z(n688) );
  CNR8X1 U959 ( .A(n688), .B(N250), .C(N274), .D(N249), .E(N270), .F(N271), 
        .G(N272), .H(N273), .Z(n689) );
  CAOR1X1 U960 ( .A(n690), .B(n689), .C(N248), .Z(N282) );
endmodule

