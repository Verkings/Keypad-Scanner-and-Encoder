
module keypad ( row, col, data, v, clock, reset );
  input [3:0] row;
  output [3:0] col;
  output [3:0] data;
  input clock, reset;
  output v;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;
  wire   [2:0] state;
  wire   [3:0] store;
  wire   [2:0] next_state;

  CFD2QX1 \state_reg[1]  ( .D(next_state[1]), .CP(clock), .CD(reset), .Q(
        state[1]) );
  CIVX2 U3 ( .A(n91), .Z(n2) );
  CIVX2 U4 ( .A(n92), .Z(n3) );
  CIVX2 U5 ( .A(n93), .Z(n4) );
  CIVX2 U6 ( .A(n94), .Z(n5) );
  CIVX2 U7 ( .A(n95), .Z(n6) );
  CIVX2 U8 ( .A(n96), .Z(n7) );
  CIVX2 U9 ( .A(n97), .Z(n8) );
  CIVX2 U10 ( .A(n98), .Z(n9) );
  CAOR1X1 U11 ( .A(col[3]), .B(n10), .C(n11), .Z(n79) );
  COND4CX1 U12 ( .A(n12), .B(n13), .C(n14), .D(n15), .Z(n10) );
  COND3X1 U13 ( .A(n16), .B(n17), .C(n18), .D(n19), .Z(n80) );
  CND2X1 U14 ( .A(col[2]), .B(n20), .Z(n19) );
  COND3X1 U15 ( .A(n21), .B(n22), .C(n23), .D(n18), .Z(n81) );
  COND4CX1 U16 ( .A(n24), .B(n25), .C(n26), .D(col[1]), .Z(n23) );
  CIVX1 U17 ( .A(n27), .Z(n26) );
  COND3X1 U18 ( .A(n21), .B(n25), .C(n18), .D(n28), .Z(n82) );
  CND2X1 U19 ( .A(col[0]), .B(n20), .Z(n28) );
  COND1XL U20 ( .A(state[0]), .B(n14), .C(n27), .Z(n20) );
  CNR2X1 U21 ( .A(n29), .B(n30), .Z(n27) );
  CAOR2X1 U22 ( .A(data[3]), .B(n31), .C(n32), .D(n33), .Z(n83) );
  CAOR2X1 U23 ( .A(data[2]), .B(n31), .C(n34), .D(n33), .Z(n84) );
  COND11X1 U24 ( .A(n35), .B(store[1]), .C(n36), .D(n37), .Z(n34) );
  COND4CX1 U25 ( .A(n38), .B(n33), .C(n39), .D(n40), .Z(n31) );
  CND2X1 U26 ( .A(n41), .B(n42), .Z(n33) );
  CNR3XL U27 ( .A(n43), .B(n13), .C(n44), .Z(n42) );
  COND1XL U28 ( .A(n45), .B(n35), .C(n46), .Z(n38) );
  CIVX1 U29 ( .A(n32), .Z(n46) );
  COND11X1 U30 ( .A(n47), .B(store[2]), .C(n48), .D(n37), .Z(n32) );
  COR3X1 U31 ( .A(n49), .B(store[3]), .C(n47), .Z(n37) );
  CND2X1 U32 ( .A(store[3]), .B(store[2]), .Z(n35) );
  COND3X1 U33 ( .A(n17), .B(n50), .C(n51), .D(n18), .Z(n85) );
  COND4CX1 U34 ( .A(n30), .B(n52), .C(n29), .D(data[1]), .Z(n51) );
  COND3X1 U35 ( .A(n17), .B(n53), .C(n54), .D(n18), .Z(n86) );
  COND1XL U36 ( .A(n29), .B(n55), .C(data[0]), .Z(n54) );
  CAOR2X1 U37 ( .A(state[0]), .B(n30), .C(n22), .D(state[1]), .Z(n55) );
  CND2IX1 U38 ( .B(n56), .A(n15), .Z(n29) );
  CANR1XL U39 ( .A(n52), .B(n57), .C(n58), .Z(n15) );
  CND3XL U40 ( .A(n59), .B(n18), .C(n60), .Z(n87) );
  COND4CX1 U41 ( .A(n61), .B(n24), .C(n62), .D(v), .Z(n60) );
  CND2X1 U42 ( .A(n12), .B(n13), .Z(n18) );
  CNR2X1 U43 ( .A(n52), .B(n63), .Z(n13) );
  COND1XL U44 ( .A(n16), .B(n24), .C(n64), .Z(n88) );
  COND4CX1 U45 ( .A(n56), .B(state[1]), .C(n65), .D(next_state[1]), .Z(n64) );
  CAOR1X1 U46 ( .A(n61), .B(n30), .C(n62), .Z(n65) );
  CNR2X1 U47 ( .A(n12), .B(n14), .Z(n30) );
  CND2X1 U48 ( .A(n66), .B(n25), .Z(n61) );
  CEOX1 U49 ( .A(state[2]), .B(n22), .Z(n66) );
  CNR2IX1 U50 ( .B(n41), .A(n43), .Z(n16) );
  CND3XL U51 ( .A(n25), .B(n63), .C(state[0]), .Z(n41) );
  COND3X1 U52 ( .A(n50), .B(n24), .C(n67), .D(n68), .Z(n89) );
  CANR2X1 U53 ( .A(next_state[2]), .B(n69), .C(n70), .D(n24), .Z(n68) );
  CIVX1 U54 ( .A(n71), .Z(n69) );
  CANR3X1 U55 ( .A(n24), .B(n52), .C(n56), .D(n62), .Z(n71) );
  CNR2IX1 U56 ( .B(n58), .A(n25), .Z(n62) );
  CNR2X1 U57 ( .A(n63), .B(n14), .Z(n56) );
  CANR11X1 U58 ( .A(state[2]), .B(n25), .C(n12), .D(n11), .Z(n67) );
  CIVX1 U59 ( .A(n59), .Z(n11) );
  CND2X1 U60 ( .A(n72), .B(n52), .Z(n59) );
  CIVX1 U61 ( .A(n44), .Z(n50) );
  CNR3XL U62 ( .A(n25), .B(state[2]), .C(n22), .Z(n44) );
  COND3X1 U63 ( .A(state[1]), .B(n73), .C(n74), .D(n75), .Z(n90) );
  CANR2X1 U64 ( .A(n14), .B(n43), .C(n39), .D(n24), .Z(n75) );
  COND1XL U65 ( .A(state[2]), .B(n52), .C(n40), .Z(n39) );
  CIVX1 U66 ( .A(n70), .Z(n40) );
  CNR3XL U67 ( .A(n63), .B(state[1]), .C(n22), .Z(n70) );
  CND2X1 U68 ( .A(n25), .B(n22), .Z(n52) );
  CIVX1 U69 ( .A(state[1]), .Z(n25) );
  CIVX1 U70 ( .A(n53), .Z(n43) );
  CND3XL U71 ( .A(n22), .B(n63), .C(state[1]), .Z(n53) );
  CANR4CX1 U73 ( .A(n58), .B(n24), .C(next_state[0]), .D(n72), .Z(n74) );
  CIVX1 U74 ( .A(n21), .Z(n72) );
  CND2X1 U75 ( .A(n12), .B(n63), .Z(n21) );
  CANR1XL U76 ( .A(n14), .B(n58), .C(n12), .Z(n73) );
  CIVX1 U77 ( .A(n17), .Z(n12) );
  CND2X1 U78 ( .A(n76), .B(n77), .Z(n17) );
  CNR2X1 U79 ( .A(n63), .B(n76), .Z(n58) );
  CIVX1 U80 ( .A(n57), .Z(n76) );
  CEOX1 U81 ( .A(n78), .B(n48), .Z(n57) );
  CIVX1 U82 ( .A(store[3]), .Z(n48) );
  CIVX1 U84 ( .A(n24), .Z(n14) );
  CND3XL U85 ( .A(n78), .B(n77), .C(store[3]), .Z(n24) );
  COND1XL U86 ( .A(n45), .B(n49), .C(n47), .Z(n77) );
  CND2X1 U87 ( .A(store[0]), .B(store[1]), .Z(n47) );
  CNR2IX1 U88 ( .B(n45), .A(n49), .Z(n78) );
  CIVX1 U89 ( .A(store[2]), .Z(n49) );
  CEOX1 U90 ( .A(store[1]), .B(n36), .Z(n45) );
  CIVX1 U91 ( .A(store[0]), .Z(n36) );
  CNR2IX1 U92 ( .B(row[0]), .A(reset), .Z(n92) );
  CNR2X1 U93 ( .A(row[0]), .B(reset), .Z(n91) );
  CNR2IX1 U94 ( .B(row[1]), .A(reset), .Z(n94) );
  CNR2X1 U95 ( .A(row[1]), .B(reset), .Z(n93) );
  CNR2IX1 U96 ( .B(row[2]), .A(reset), .Z(n96) );
  CNR2X1 U97 ( .A(row[2]), .B(reset), .Z(n95) );
  CNR2IX1 U98 ( .B(row[3]), .A(reset), .Z(n98) );
  CNR2X1 U99 ( .A(row[3]), .B(reset), .Z(n97) );
  CFD3QXL \store_reg[3]  ( .D(row[3]), .CP(clock), .CD(n8), .SD(n9), .Q(
        store[3]) );
  CFD3QXL \store_reg[2]  ( .D(row[2]), .CP(clock), .CD(n6), .SD(n7), .Q(
        store[2]) );
  CFD3QXL \store_reg[1]  ( .D(row[1]), .CP(clock), .CD(n4), .SD(n5), .Q(
        store[1]) );
  CFD3QXL \store_reg[0]  ( .D(row[0]), .CP(clock), .CD(n2), .SD(n3), .Q(
        store[0]) );
  CFD2XL \state_reg[2]  ( .D(next_state[2]), .CP(clock), .CD(reset), .Q(
        state[2]), .QN(n63) );
  CFD1QXL \data_reg[3]  ( .D(n83), .CP(clock), .Q(data[3]) );
  CFD1QXL \data_reg[2]  ( .D(n84), .CP(clock), .Q(data[2]) );
  CFD1QXL v_reg ( .D(n87), .CP(clock), .Q(v) );
  CFD1QXL \col_reg[3]  ( .D(n79), .CP(clock), .Q(col[3]) );
  CFD1QXL \next_state_reg[0]  ( .D(n90), .CP(clock), .Q(next_state[0]) );
  CFD1QXL \next_state_reg[1]  ( .D(n88), .CP(clock), .Q(next_state[1]) );
  CFD1QXL \data_reg[1]  ( .D(n85), .CP(clock), .Q(data[1]) );
  CFD1QXL \data_reg[0]  ( .D(n86), .CP(clock), .Q(data[0]) );
  CFD1QXL \col_reg[1]  ( .D(n81), .CP(clock), .Q(col[1]) );
  CFD1QXL \next_state_reg[2]  ( .D(n89), .CP(clock), .Q(next_state[2]) );
  CFD1QXL \col_reg[2]  ( .D(n80), .CP(clock), .Q(col[2]) );
  CFD1QXL \col_reg[0]  ( .D(n82), .CP(clock), .Q(col[0]) );
  CFD2XL \state_reg[0]  ( .D(next_state[0]), .CP(clock), .CD(reset), .Q(
        state[0]), .QN(n22) );
endmodule


module controller ( v, clock, reset, full, empty, read, valid, wr_enable, 
        rd_enable );
  input v, clock, reset, full, empty, read;
  output valid, wr_enable, rd_enable;
  wire   N19, N20, N21, n1;
  assign N20 = v;

  CFD2QX1 wr_enable_reg ( .D(N20), .CP(clock), .CD(reset), .Q(wr_enable) );
  CFD4QXL valid_reg ( .D(N21), .CP(clock), .SD(reset), .Q(valid) );
  CNR2X1 U3 ( .A(read), .B(n1), .Z(N21) );
  CNR2IX1 U4 ( .B(read), .A(n1), .Z(N19) );
  CNR2IX1 U5 ( .B(empty), .A(N20), .Z(n1) );
  CFD2QX2 rd_enable_reg ( .D(N19), .CP(clock), .CD(reset), .Q(rd_enable) );
endmodule


module fifo_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B_not[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59;
  wire   [32:0] carry;

  CENXL U1 ( .A(A[19]), .B(carry[19]), .Z(DIFF[19]) );
  CENXL U2 ( .A(A[5]), .B(carry[5]), .Z(DIFF[5]) );
  CENXL U3 ( .A(A[20]), .B(carry[20]), .Z(DIFF[20]) );
  CENXL U4 ( .A(A[25]), .B(carry[25]), .Z(DIFF[25]) );
  CENXL U5 ( .A(A[10]), .B(carry[10]), .Z(DIFF[10]) );
  CENXL U6 ( .A(A[26]), .B(carry[26]), .Z(DIFF[26]) );
  CENXL U7 ( .A(A[15]), .B(carry[15]), .Z(DIFF[15]) );
  CENXL U8 ( .A(A[12]), .B(carry[12]), .Z(DIFF[12]) );
  CIVX2 U9 ( .A(carry[3]), .Z(n1) );
  CIVDXL U10 ( .A(carry[3]), .Z1(n2) );
  CNR2IX1 U11 ( .B(n45), .A(carry[30]), .Z(n4) );
  CENX1 U12 ( .A(A[3]), .B(n2), .Z(DIFF[3]) );
  CND2IX2 U13 ( .B(A[27]), .A(n38), .Z(carry[28]) );
  CENX1 U14 ( .A(A[28]), .B(carry[28]), .Z(DIFF[28]) );
  CENX1 U15 ( .A(A[30]), .B(carry[30]), .Z(DIFF[30]) );
  CENX1 U16 ( .A(n3), .B(n4), .Z(DIFF[31]) );
  CIVX20 U17 ( .A(A[31]), .Z(n3) );
  CENX1 U18 ( .A(A[29]), .B(carry[29]), .Z(DIFF[29]) );
  CND2IX2 U19 ( .B(A[17]), .A(n18), .Z(carry[18]) );
  CIVX2 U20 ( .A(B[0]), .Z(\B_not[0] ) );
  CENXL U21 ( .A(\B_not[0] ), .B(A[0]), .Z(DIFF[0]) );
  CND2IX2 U22 ( .B(A[13]), .A(n11), .Z(carry[14]) );
  CND2IX2 U23 ( .B(A[21]), .A(n27), .Z(carry[22]) );
  CENXL U24 ( .A(A[24]), .B(carry[24]), .Z(DIFF[24]) );
  CENXL U25 ( .A(A[2]), .B(carry[2]), .Z(DIFF[2]) );
  CENXL U26 ( .A(A[9]), .B(carry[9]), .Z(DIFF[9]) );
  CENXL U27 ( .A(A[18]), .B(carry[18]), .Z(DIFF[18]) );
  CENXL U28 ( .A(A[8]), .B(carry[8]), .Z(DIFF[8]) );
  CENXL U29 ( .A(A[16]), .B(carry[16]), .Z(DIFF[16]) );
  CENXL U30 ( .A(A[1]), .B(carry[1]), .Z(DIFF[1]) );
  CENXL U31 ( .A(A[7]), .B(carry[7]), .Z(DIFF[7]) );
  CENXL U32 ( .A(A[6]), .B(carry[6]), .Z(DIFF[6]) );
  CENXL U33 ( .A(A[21]), .B(carry[21]), .Z(DIFF[21]) );
  CENXL U34 ( .A(A[22]), .B(carry[22]), .Z(DIFF[22]) );
  CENXL U35 ( .A(A[13]), .B(carry[13]), .Z(DIFF[13]) );
  CENXL U36 ( .A(A[14]), .B(carry[14]), .Z(DIFF[14]) );
  CENXL U37 ( .A(A[4]), .B(carry[4]), .Z(DIFF[4]) );
  CENXL U38 ( .A(A[17]), .B(carry[17]), .Z(DIFF[17]) );
  CENXL U39 ( .A(A[23]), .B(carry[23]), .Z(DIFF[23]) );
  CENXL U40 ( .A(A[11]), .B(carry[11]), .Z(DIFF[11]) );
  CND2X2 U41 ( .A(n5), .B(n6), .Z(carry[11]) );
  CIVX2 U42 ( .A(A[10]), .Z(n5) );
  CIVX2 U43 ( .A(carry[10]), .Z(n6) );
  CND2X2 U44 ( .A(n7), .B(n8), .Z(carry[12]) );
  CIVX2 U45 ( .A(A[11]), .Z(n7) );
  CIVX2 U46 ( .A(carry[11]), .Z(n8) );
  CND2X2 U47 ( .A(n9), .B(n10), .Z(carry[13]) );
  CIVX2 U48 ( .A(A[12]), .Z(n9) );
  CIVX2 U49 ( .A(carry[12]), .Z(n10) );
  CIVX2 U50 ( .A(carry[13]), .Z(n11) );
  CND2X2 U51 ( .A(n12), .B(n13), .Z(carry[15]) );
  CIVX2 U52 ( .A(A[14]), .Z(n12) );
  CIVX2 U53 ( .A(carry[14]), .Z(n13) );
  CND2X2 U54 ( .A(n14), .B(n15), .Z(carry[16]) );
  CIVX2 U55 ( .A(A[15]), .Z(n14) );
  CIVX2 U56 ( .A(carry[15]), .Z(n15) );
  CND2X2 U57 ( .A(n16), .B(n17), .Z(carry[17]) );
  CIVX2 U58 ( .A(A[16]), .Z(n16) );
  CIVX2 U59 ( .A(carry[16]), .Z(n17) );
  CIVX2 U60 ( .A(carry[17]), .Z(n18) );
  CND2X2 U61 ( .A(n19), .B(n20), .Z(carry[19]) );
  CIVX2 U62 ( .A(A[18]), .Z(n19) );
  CIVX2 U63 ( .A(carry[18]), .Z(n20) );
  CND2X2 U64 ( .A(n21), .B(n22), .Z(carry[20]) );
  CIVX2 U65 ( .A(A[19]), .Z(n21) );
  CIVX2 U66 ( .A(carry[19]), .Z(n22) );
  CND2X2 U67 ( .A(n24), .B(n23), .Z(carry[2]) );
  CIVX2 U68 ( .A(A[1]), .Z(n23) );
  CIVX2 U69 ( .A(carry[1]), .Z(n24) );
  CND2X2 U70 ( .A(n25), .B(n26), .Z(carry[21]) );
  CIVX2 U71 ( .A(A[20]), .Z(n25) );
  CIVX2 U72 ( .A(carry[20]), .Z(n26) );
  CIVX2 U73 ( .A(carry[21]), .Z(n27) );
  CND2X2 U74 ( .A(n28), .B(n29), .Z(carry[23]) );
  CIVX2 U75 ( .A(A[22]), .Z(n28) );
  CIVX2 U76 ( .A(carry[22]), .Z(n29) );
  CND2X2 U77 ( .A(n30), .B(n31), .Z(carry[24]) );
  CIVX2 U78 ( .A(A[23]), .Z(n30) );
  CIVX2 U79 ( .A(carry[23]), .Z(n31) );
  CND2X2 U80 ( .A(n32), .B(n33), .Z(carry[25]) );
  CIVX2 U81 ( .A(A[24]), .Z(n32) );
  CIVX2 U82 ( .A(carry[24]), .Z(n33) );
  CND2X2 U83 ( .A(n34), .B(n35), .Z(carry[26]) );
  CIVX2 U84 ( .A(A[25]), .Z(n34) );
  CIVX2 U85 ( .A(carry[25]), .Z(n35) );
  CND2X2 U86 ( .A(n36), .B(n37), .Z(carry[27]) );
  CIVX2 U87 ( .A(A[26]), .Z(n36) );
  CIVX2 U88 ( .A(carry[26]), .Z(n37) );
  CENX2 U89 ( .A(A[27]), .B(carry[27]), .Z(DIFF[27]) );
  CIVX2 U90 ( .A(carry[27]), .Z(n38) );
  CND2X2 U91 ( .A(n40), .B(n39), .Z(carry[29]) );
  CIVX2 U92 ( .A(A[28]), .Z(n39) );
  CIVX2 U93 ( .A(carry[28]), .Z(n40) );
  CND2X2 U94 ( .A(n41), .B(n42), .Z(carry[30]) );
  CIVX2 U95 ( .A(A[29]), .Z(n41) );
  CIVX2 U96 ( .A(carry[29]), .Z(n42) );
  CND2X2 U97 ( .A(n44), .B(n43), .Z(carry[3]) );
  CIVX2 U98 ( .A(A[2]), .Z(n43) );
  CIVX2 U99 ( .A(carry[2]), .Z(n44) );
  CIVX2 U100 ( .A(A[30]), .Z(n45) );
  CND2X2 U101 ( .A(n1), .B(n46), .Z(carry[4]) );
  CIVX2 U102 ( .A(A[3]), .Z(n46) );
  CND2X2 U103 ( .A(n47), .B(n48), .Z(carry[5]) );
  CIVX2 U104 ( .A(A[4]), .Z(n47) );
  CIVX2 U105 ( .A(carry[4]), .Z(n48) );
  CND2X2 U106 ( .A(n49), .B(n50), .Z(carry[6]) );
  CIVX2 U107 ( .A(A[5]), .Z(n49) );
  CIVX2 U108 ( .A(carry[5]), .Z(n50) );
  CND2X2 U109 ( .A(n52), .B(n51), .Z(carry[7]) );
  CIVX2 U110 ( .A(A[6]), .Z(n51) );
  CIVX2 U111 ( .A(carry[6]), .Z(n52) );
  CND2X2 U112 ( .A(n54), .B(n53), .Z(carry[8]) );
  CIVX2 U113 ( .A(A[7]), .Z(n53) );
  CIVX2 U114 ( .A(carry[7]), .Z(n54) );
  CND2X2 U115 ( .A(n56), .B(n55), .Z(carry[9]) );
  CIVX2 U116 ( .A(A[8]), .Z(n55) );
  CIVX2 U117 ( .A(carry[8]), .Z(n56) );
  CND2X2 U118 ( .A(n57), .B(n58), .Z(carry[10]) );
  CIVX2 U119 ( .A(A[9]), .Z(n57) );
  CIVX2 U120 ( .A(carry[9]), .Z(n58) );
  CND2X2 U121 ( .A(B[0]), .B(n59), .Z(carry[1]) );
  CIVX2 U122 ( .A(A[0]), .Z(n59) );
endmodule


module fifo_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91;
  assign n49 = A[11];
  assign n58 = A[9];
  assign n65 = A[7];
  assign n73 = A[5];
  assign n77 = A[4];
  assign n82 = A[3];
  assign n85 = A[2];
  assign n89 = A[1];
  assign n91 = A[0];

  CEOX2 U1 ( .A(A[31]), .B(n1), .Z(SUM[31]) );
  CHA1X1 U2 ( .A(A[30]), .B(n2), .CO(n1), .S(SUM[30]) );
  CHA1X1 U3 ( .A(A[29]), .B(n3), .CO(n2), .S(SUM[29]) );
  CHA1X1 U4 ( .A(A[28]), .B(n4), .CO(n3), .S(SUM[28]) );
  CHA1X1 U5 ( .A(A[27]), .B(n5), .CO(n4), .S(SUM[27]) );
  CHA1X1 U6 ( .A(A[26]), .B(n6), .CO(n5), .S(SUM[26]) );
  CHA1X1 U7 ( .A(A[25]), .B(n7), .CO(n6), .S(SUM[25]) );
  CHA1X1 U8 ( .A(A[24]), .B(n8), .CO(n7), .S(SUM[24]) );
  CEOX2 U9 ( .A(n11), .B(n12), .Z(SUM[23]) );
  CNR2X2 U10 ( .A(n9), .B(n52), .Z(n8) );
  CND2X2 U11 ( .A(n26), .B(n10), .Z(n9) );
  CNR2X2 U12 ( .A(n14), .B(n11), .Z(n10) );
  CENX2 U14 ( .A(n17), .B(n16), .Z(SUM[22]) );
  CND2X2 U15 ( .A(n24), .B(n13), .Z(n12) );
  CND2X2 U17 ( .A(n15), .B(n20), .Z(n14) );
  CNR2X2 U18 ( .A(n16), .B(n18), .Z(n15) );
  CEOX2 U20 ( .A(n18), .B(n19), .Z(SUM[21]) );
  CNR2X2 U21 ( .A(n19), .B(n18), .Z(n17) );
  CENX2 U23 ( .A(n22), .B(n21), .Z(SUM[20]) );
  CND2X2 U24 ( .A(n24), .B(n20), .Z(n19) );
  CNR2X2 U25 ( .A(n21), .B(n23), .Z(n20) );
  CENX2 U27 ( .A(n24), .B(n23), .Z(SUM[19]) );
  CNR2X2 U28 ( .A(n25), .B(n23), .Z(n22) );
  CENX2 U30 ( .A(n30), .B(n29), .Z(SUM[18]) );
  CND2X2 U32 ( .A(n51), .B(n26), .Z(n25) );
  CNR2X2 U33 ( .A(n40), .B(n27), .Z(n26) );
  CND2X2 U34 ( .A(n33), .B(n28), .Z(n27) );
  CNR2X2 U35 ( .A(n31), .B(n29), .Z(n28) );
  CEOX2 U37 ( .A(n31), .B(n32), .Z(SUM[17]) );
  CNR2X2 U38 ( .A(n32), .B(n31), .Z(n30) );
  CENX2 U40 ( .A(n35), .B(n34), .Z(SUM[16]) );
  CND2X2 U41 ( .A(n37), .B(n33), .Z(n32) );
  CNR2X2 U42 ( .A(n34), .B(n36), .Z(n33) );
  CENX2 U44 ( .A(n37), .B(n36), .Z(SUM[15]) );
  CNR2X2 U45 ( .A(n38), .B(n36), .Z(n35) );
  CENX2 U47 ( .A(n43), .B(n42), .Z(SUM[14]) );
  CND2X2 U49 ( .A(n51), .B(n39), .Z(n38) );
  CND2X2 U51 ( .A(n41), .B(n46), .Z(n40) );
  CNR2X2 U52 ( .A(n42), .B(n44), .Z(n41) );
  CEOX2 U54 ( .A(n44), .B(n45), .Z(SUM[13]) );
  CNR2X2 U55 ( .A(n45), .B(n44), .Z(n43) );
  CEOX2 U57 ( .A(n47), .B(n48), .Z(SUM[12]) );
  CND2X2 U58 ( .A(n51), .B(n46), .Z(n45) );
  CNR2X2 U59 ( .A(n47), .B(n50), .Z(n46) );
  CENX2 U61 ( .A(n51), .B(n50), .Z(SUM[11]) );
  CND2X2 U62 ( .A(n51), .B(n49), .Z(n48) );
  CEOX2 U65 ( .A(n56), .B(n57), .Z(SUM[10]) );
  CND2X2 U67 ( .A(n53), .B(n80), .Z(n52) );
  CNR2X2 U68 ( .A(n54), .B(n69), .Z(n53) );
  CND2X2 U69 ( .A(n62), .B(n55), .Z(n54) );
  CNR2X2 U70 ( .A(n56), .B(n59), .Z(n55) );
  CENX2 U72 ( .A(n60), .B(n59), .Z(SUM[9]) );
  CND2X2 U73 ( .A(n60), .B(n58), .Z(n57) );
  CEOX2 U76 ( .A(n63), .B(n64), .Z(SUM[8]) );
  CNR2X2 U77 ( .A(n67), .B(n61), .Z(n60) );
  CNR2X2 U79 ( .A(n63), .B(n66), .Z(n62) );
  CEOX2 U81 ( .A(n66), .B(n67), .Z(SUM[7]) );
  CND2X2 U82 ( .A(n68), .B(n65), .Z(n64) );
  CEOX2 U85 ( .A(n71), .B(n72), .Z(SUM[6]) );
  CNR2X2 U87 ( .A(n79), .B(n69), .Z(n68) );
  CND2X2 U88 ( .A(n70), .B(n77), .Z(n69) );
  CNR2X2 U89 ( .A(n71), .B(n74), .Z(n70) );
  CENX2 U91 ( .A(n75), .B(n74), .Z(SUM[5]) );
  CND2X2 U92 ( .A(n75), .B(n73), .Z(n72) );
  CEOX2 U95 ( .A(n78), .B(n79), .Z(SUM[4]) );
  CNR2X2 U96 ( .A(n79), .B(n78), .Z(n75) );
  CEOX2 U100 ( .A(n83), .B(n84), .Z(SUM[3]) );
  CNR2X2 U102 ( .A(n81), .B(n88), .Z(n80) );
  CND2X2 U103 ( .A(n85), .B(n82), .Z(n81) );
  CENX2 U106 ( .A(n86), .B(n87), .Z(SUM[2]) );
  CND2X2 U107 ( .A(n87), .B(n85), .Z(n84) );
  CENX2 U110 ( .A(n90), .B(n91), .Z(SUM[1]) );
  CND2X2 U112 ( .A(n91), .B(n89), .Z(n88) );
  CIVX2 U119 ( .A(n89), .Z(n90) );
  CIVX2 U120 ( .A(n88), .Z(n87) );
  CIVX2 U121 ( .A(n85), .Z(n86) );
  CIVX2 U122 ( .A(n82), .Z(n83) );
  CIVX2 U123 ( .A(n80), .Z(n79) );
  CIVX2 U124 ( .A(n77), .Z(n78) );
  CIVX2 U125 ( .A(n73), .Z(n74) );
  CIVX2 U126 ( .A(A[6]), .Z(n71) );
  CIVX2 U127 ( .A(n68), .Z(n67) );
  CIVX2 U128 ( .A(n65), .Z(n66) );
  CIVX2 U129 ( .A(A[8]), .Z(n63) );
  CIVX2 U130 ( .A(n62), .Z(n61) );
  CIVX2 U131 ( .A(n58), .Z(n59) );
  CIVX2 U132 ( .A(A[10]), .Z(n56) );
  CIVX2 U133 ( .A(n52), .Z(n51) );
  CIVX2 U134 ( .A(n49), .Z(n50) );
  CIVX2 U135 ( .A(A[12]), .Z(n47) );
  CIVX2 U136 ( .A(A[13]), .Z(n44) );
  CIVX2 U137 ( .A(A[14]), .Z(n42) );
  CIVX2 U138 ( .A(n40), .Z(n39) );
  CIVX2 U139 ( .A(n38), .Z(n37) );
  CIVX2 U140 ( .A(A[15]), .Z(n36) );
  CIVX2 U141 ( .A(A[16]), .Z(n34) );
  CIVX2 U142 ( .A(A[17]), .Z(n31) );
  CIVX2 U143 ( .A(A[18]), .Z(n29) );
  CIVX2 U144 ( .A(n25), .Z(n24) );
  CIVX2 U145 ( .A(A[19]), .Z(n23) );
  CIVX2 U146 ( .A(A[20]), .Z(n21) );
  CIVX2 U147 ( .A(A[21]), .Z(n18) );
  CIVX2 U148 ( .A(A[22]), .Z(n16) );
  CIVX2 U149 ( .A(n14), .Z(n13) );
  CIVX2 U150 ( .A(A[23]), .Z(n11) );
  CIVX2 U151 ( .A(n91), .Z(SUM[0]) );
endmodule


module fifo ( code, full, empty, data, rd_enable, wr_enable, reset, clock );
  output [3:0] code;
  input [3:0] data;
  input rd_enable, wr_enable, reset, clock;
  output full, empty;
  wire   N50, \memory[31][3] , \memory[31][2] , \memory[31][1] ,
         \memory[31][0] , \memory[30][3] , \memory[30][2] , \memory[30][1] ,
         \memory[30][0] , \memory[29][3] , \memory[29][2] , \memory[29][1] ,
         \memory[29][0] , \memory[28][3] , \memory[28][2] , \memory[28][1] ,
         \memory[28][0] , \memory[27][3] , \memory[27][2] , \memory[27][1] ,
         \memory[27][0] , \memory[26][3] , \memory[26][2] , \memory[26][1] ,
         \memory[26][0] , \memory[25][3] , \memory[25][2] , \memory[25][1] ,
         \memory[25][0] , \memory[24][3] , \memory[24][2] , \memory[24][1] ,
         \memory[24][0] , \memory[23][3] , \memory[23][2] , \memory[23][1] ,
         \memory[23][0] , \memory[22][3] , \memory[22][2] , \memory[22][1] ,
         \memory[22][0] , \memory[21][3] , \memory[21][2] , \memory[21][1] ,
         \memory[21][0] , \memory[20][3] , \memory[20][2] , \memory[20][1] ,
         \memory[20][0] , \memory[19][3] , \memory[19][2] , \memory[19][1] ,
         \memory[19][0] , \memory[18][3] , \memory[18][2] , \memory[18][1] ,
         \memory[18][0] , \memory[17][3] , \memory[17][2] , \memory[17][1] ,
         \memory[17][0] , \memory[16][3] , \memory[16][2] , \memory[16][1] ,
         \memory[16][0] , \memory[15][3] , \memory[15][2] , \memory[15][1] ,
         \memory[15][0] , \memory[14][3] , \memory[14][2] , \memory[14][1] ,
         \memory[14][0] , \memory[13][3] , \memory[13][2] , \memory[13][1] ,
         \memory[13][0] , \memory[12][3] , \memory[12][2] , \memory[12][1] ,
         \memory[12][0] , \memory[11][3] , \memory[11][2] , \memory[11][1] ,
         \memory[11][0] , \memory[10][3] , \memory[10][2] , \memory[10][1] ,
         \memory[10][0] , \memory[9][3] , \memory[9][2] , \memory[9][1] ,
         \memory[9][0] , \memory[8][3] , \memory[8][2] , \memory[8][1] ,
         \memory[8][0] , \memory[7][3] , \memory[7][2] , \memory[7][1] ,
         \memory[7][0] , \memory[6][3] , \memory[6][2] , \memory[6][1] ,
         \memory[6][0] , \memory[5][3] , \memory[5][2] , \memory[5][1] ,
         \memory[5][0] , \memory[4][3] , \memory[4][2] , \memory[4][1] ,
         \memory[4][0] , \memory[3][3] , \memory[3][2] , \memory[3][1] ,
         \memory[3][0] , \memory[2][3] , \memory[2][2] , \memory[2][1] ,
         \memory[2][0] , \memory[0][3] , \memory[0][2] , \memory[0][1] ,
         \memory[0][0] , N61, N63, N65, N67, N69, N71, N73, N75, N77, N79, N81,
         N83, N85, N87, N89, N91, N93, N95, N97, N99, N101, N103, N105, N107,
         N109, N111, N113, N115, N117, N119, N121, N123, N248, N249, N250,
         N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261,
         N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272,
         N273, N274, N275, N276, N277, N278, N279, N282, N563, N564, N565,
         N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576,
         N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587,
         N588, N589, N590, N591, N592, N593, N594, N1652, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n14, n15, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852;
  wire   [31:0] counter;

  CFD2QX1 \counter_reg[0]  ( .D(n790), .CP(clock), .CD(reset), .Q(counter[0])
         );
  CFD2QX1 \counter_reg[31]  ( .D(n789), .CP(clock), .CD(reset), .Q(counter[31]) );
  CFD2QX1 \counter_reg[1]  ( .D(n788), .CP(clock), .CD(reset), .Q(counter[1])
         );
  CFD2QX1 \counter_reg[30]  ( .D(n759), .CP(clock), .CD(reset), .Q(counter[30]) );
  CFD2QX1 \counter_reg[2]  ( .D(n787), .CP(clock), .CD(reset), .Q(counter[2])
         );
  CFD2QX1 \counter_reg[3]  ( .D(n786), .CP(clock), .CD(reset), .Q(counter[3])
         );
  CFD2QX1 \counter_reg[4]  ( .D(n785), .CP(clock), .CD(reset), .Q(counter[4])
         );
  CFD2QX1 \counter_reg[5]  ( .D(n784), .CP(clock), .CD(reset), .Q(counter[5])
         );
  CFD2QX1 \counter_reg[6]  ( .D(n783), .CP(clock), .CD(reset), .Q(counter[6])
         );
  CFD2QX1 \counter_reg[7]  ( .D(n782), .CP(clock), .CD(reset), .Q(counter[7])
         );
  CFD2QX1 \counter_reg[8]  ( .D(n781), .CP(clock), .CD(reset), .Q(counter[8])
         );
  CFD2QX1 \counter_reg[9]  ( .D(n780), .CP(clock), .CD(reset), .Q(counter[9])
         );
  CFD2QX1 \counter_reg[10]  ( .D(n779), .CP(clock), .CD(reset), .Q(counter[10]) );
  CFD2QX1 \counter_reg[11]  ( .D(n778), .CP(clock), .CD(reset), .Q(counter[11]) );
  CFD2QX1 \counter_reg[12]  ( .D(n777), .CP(clock), .CD(reset), .Q(counter[12]) );
  CFD2QX1 \counter_reg[13]  ( .D(n776), .CP(clock), .CD(reset), .Q(counter[13]) );
  CFD2QX1 \counter_reg[14]  ( .D(n775), .CP(clock), .CD(reset), .Q(counter[14]) );
  CFD2QX1 \counter_reg[15]  ( .D(n774), .CP(clock), .CD(reset), .Q(counter[15]) );
  CFD2QX1 \counter_reg[16]  ( .D(n773), .CP(clock), .CD(reset), .Q(counter[16]) );
  CFD2QX1 \counter_reg[17]  ( .D(n772), .CP(clock), .CD(reset), .Q(counter[17]) );
  CFD2QX1 \counter_reg[18]  ( .D(n771), .CP(clock), .CD(reset), .Q(counter[18]) );
  CFD2QX1 \counter_reg[19]  ( .D(n770), .CP(clock), .CD(reset), .Q(counter[19]) );
  CFD2QX1 \counter_reg[20]  ( .D(n769), .CP(clock), .CD(reset), .Q(counter[20]) );
  CFD2QX1 \counter_reg[21]  ( .D(n768), .CP(clock), .CD(reset), .Q(counter[21]) );
  CFD2QX1 \counter_reg[22]  ( .D(n767), .CP(clock), .CD(reset), .Q(counter[22]) );
  CFD2QX1 \counter_reg[23]  ( .D(n766), .CP(clock), .CD(reset), .Q(counter[23]) );
  CFD2QX1 \counter_reg[24]  ( .D(n765), .CP(clock), .CD(reset), .Q(counter[24]) );
  CFD2QX1 \counter_reg[25]  ( .D(n764), .CP(clock), .CD(reset), .Q(counter[25]) );
  CFD2QX1 \counter_reg[26]  ( .D(n763), .CP(clock), .CD(reset), .Q(counter[26]) );
  CFD2QX1 \counter_reg[27]  ( .D(n762), .CP(clock), .CD(reset), .Q(counter[27]) );
  CFD2QX1 \counter_reg[28]  ( .D(n761), .CP(clock), .CD(reset), .Q(counter[28]) );
  CFD2QX1 \counter_reg[29]  ( .D(n760), .CP(clock), .CD(reset), .Q(counter[29]) );
  CFD4QXL empty_reg ( .D(n626), .CP(clock), .SD(reset), .Q(empty) );
  CFD2QX1 full_reg ( .D(n625), .CP(clock), .CD(reset), .Q(full) );
  CAOR2X1 U3 ( .A(full), .B(n16), .C(n17), .D(n18), .Z(n625) );
  CIVX1 U10 ( .A(n20), .Z(n19) );
  CANR1XL U11 ( .A(n21), .B(n22), .C(N1652), .Z(n20) );
  COND1XL U12 ( .A(n23), .B(n24), .C(n25), .Z(n627) );
  CANR2X1 U13 ( .A(\memory[31][3] ), .B(n26), .C(n27), .D(n28), .Z(n25) );
  COND1XL U14 ( .A(n23), .B(n29), .C(n30), .Z(n628) );
  CANR2X1 U15 ( .A(\memory[31][2] ), .B(n26), .C(n31), .D(n28), .Z(n30) );
  COND1XL U16 ( .A(n23), .B(n32), .C(n33), .Z(n629) );
  CANR2X1 U17 ( .A(\memory[31][1] ), .B(n26), .C(n34), .D(n28), .Z(n33) );
  COND1XL U18 ( .A(n23), .B(n35), .C(n36), .Z(n630) );
  CANR2X1 U19 ( .A(\memory[31][0] ), .B(n26), .C(n37), .D(n28), .Z(n36) );
  CNR2IX1 U20 ( .B(n23), .A(n38), .Z(n28) );
  COAN1X1 U21 ( .A(n38), .B(n21), .C(n23), .Z(n26) );
  COND1XL U22 ( .A(n39), .B(n38), .C(n16), .Z(n23) );
  CND2X1 U23 ( .A(n40), .B(n41), .Z(n38) );
  COND1XL U24 ( .A(n42), .B(n43), .C(n44), .Z(n631) );
  COND4CX1 U25 ( .A(n45), .B(\memory[31][3] ), .C(n46), .D(n42), .Z(n44) );
  COND2X1 U26 ( .A(n793), .B(n24), .C(n48), .D(n49), .Z(n46) );
  COND1XL U27 ( .A(n42), .B(n50), .C(n51), .Z(n632) );
  COND4CX1 U28 ( .A(n45), .B(\memory[31][2] ), .C(n52), .D(n42), .Z(n51) );
  COND2X1 U29 ( .A(n793), .B(n29), .C(n53), .D(n49), .Z(n52) );
  COND1XL U30 ( .A(n42), .B(n54), .C(n55), .Z(n633) );
  COND4CX1 U31 ( .A(n45), .B(\memory[31][1] ), .C(n56), .D(n42), .Z(n55) );
  COND2X1 U32 ( .A(n793), .B(n32), .C(n57), .D(n49), .Z(n56) );
  COND1XL U33 ( .A(n42), .B(n58), .C(n59), .Z(n634) );
  COND4CX1 U34 ( .A(n45), .B(\memory[31][0] ), .C(n60), .D(n42), .Z(n59) );
  COND2X1 U35 ( .A(n793), .B(n35), .C(n61), .D(n49), .Z(n60) );
  CANR1XL U36 ( .A(n49), .B(N282), .C(n62), .Z(n47) );
  COND1XL U37 ( .A(n39), .B(n49), .C(n16), .Z(n42) );
  CND2X1 U38 ( .A(n63), .B(n40), .Z(n49) );
  COND1XL U39 ( .A(n64), .B(n65), .C(n66), .Z(n635) );
  COND4CX1 U40 ( .A(n45), .B(\memory[30][3] ), .C(n67), .D(n64), .Z(n66) );
  COND2X1 U41 ( .A(n795), .B(n43), .C(n48), .D(n69), .Z(n67) );
  COND1XL U42 ( .A(n64), .B(n70), .C(n71), .Z(n636) );
  COND4CX1 U43 ( .A(n45), .B(\memory[30][2] ), .C(n72), .D(n64), .Z(n71) );
  COND2X1 U44 ( .A(n795), .B(n50), .C(n53), .D(n69), .Z(n72) );
  COND1XL U45 ( .A(n64), .B(n73), .C(n74), .Z(n637) );
  COND4CX1 U46 ( .A(n45), .B(\memory[30][1] ), .C(n75), .D(n64), .Z(n74) );
  COND2X1 U47 ( .A(n795), .B(n54), .C(n57), .D(n69), .Z(n75) );
  COND1XL U48 ( .A(n64), .B(n76), .C(n77), .Z(n638) );
  COND4CX1 U49 ( .A(n45), .B(\memory[30][0] ), .C(n78), .D(n64), .Z(n77) );
  COND2X1 U50 ( .A(n795), .B(n58), .C(n61), .D(n69), .Z(n78) );
  CANR1XL U51 ( .A(n69), .B(N282), .C(n62), .Z(n68) );
  COND1XL U52 ( .A(n39), .B(n69), .C(n16), .Z(n64) );
  CND2X1 U53 ( .A(n79), .B(n40), .Z(n69) );
  COND1XL U54 ( .A(n80), .B(n81), .C(n82), .Z(n639) );
  COND4CX1 U55 ( .A(\memory[29][3] ), .B(n45), .C(n83), .D(n80), .Z(n82) );
  COND2X1 U56 ( .A(n797), .B(n65), .C(n48), .D(n85), .Z(n83) );
  COND1XL U57 ( .A(n80), .B(n86), .C(n87), .Z(n640) );
  COND4CX1 U58 ( .A(\memory[29][2] ), .B(n45), .C(n88), .D(n80), .Z(n87) );
  COND2X1 U59 ( .A(n797), .B(n70), .C(n53), .D(n85), .Z(n88) );
  COND1XL U60 ( .A(n80), .B(n89), .C(n90), .Z(n641) );
  COND4CX1 U61 ( .A(\memory[29][1] ), .B(n45), .C(n91), .D(n80), .Z(n90) );
  COND2X1 U62 ( .A(n797), .B(n73), .C(n57), .D(n85), .Z(n91) );
  COND1XL U63 ( .A(n80), .B(n92), .C(n93), .Z(n642) );
  COND4CX1 U64 ( .A(\memory[29][0] ), .B(n45), .C(n94), .D(n80), .Z(n93) );
  COND2X1 U65 ( .A(n797), .B(n76), .C(n61), .D(n85), .Z(n94) );
  CANR1XL U66 ( .A(n85), .B(N282), .C(n62), .Z(n84) );
  COND1XL U67 ( .A(n39), .B(n85), .C(n16), .Z(n80) );
  CND2X1 U68 ( .A(n95), .B(n40), .Z(n85) );
  COND1XL U69 ( .A(n96), .B(n97), .C(n98), .Z(n643) );
  COND4CX1 U70 ( .A(\memory[28][3] ), .B(n45), .C(n99), .D(n96), .Z(n98) );
  COND2X1 U71 ( .A(n799), .B(n81), .C(n48), .D(n101), .Z(n99) );
  COND1XL U72 ( .A(n96), .B(n102), .C(n103), .Z(n644) );
  COND4CX1 U73 ( .A(\memory[28][2] ), .B(n45), .C(n104), .D(n96), .Z(n103) );
  COND2X1 U74 ( .A(n799), .B(n86), .C(n53), .D(n101), .Z(n104) );
  COND1XL U75 ( .A(n96), .B(n105), .C(n106), .Z(n645) );
  COND4CX1 U76 ( .A(\memory[28][1] ), .B(n45), .C(n107), .D(n96), .Z(n106) );
  COND2X1 U77 ( .A(n799), .B(n89), .C(n57), .D(n101), .Z(n107) );
  COND1XL U78 ( .A(n96), .B(n108), .C(n109), .Z(n646) );
  COND4CX1 U79 ( .A(\memory[28][0] ), .B(n45), .C(n110), .D(n96), .Z(n109) );
  COND2X1 U80 ( .A(n799), .B(n92), .C(n61), .D(n101), .Z(n110) );
  CANR1XL U81 ( .A(n101), .B(N282), .C(n62), .Z(n100) );
  COND1XL U82 ( .A(n39), .B(n101), .C(n16), .Z(n96) );
  CND2X1 U83 ( .A(n111), .B(n40), .Z(n101) );
  COND1XL U84 ( .A(n112), .B(n113), .C(n114), .Z(n647) );
  COND4CX1 U85 ( .A(\memory[27][3] ), .B(n45), .C(n115), .D(n112), .Z(n114) );
  COND2X1 U86 ( .A(n801), .B(n97), .C(n48), .D(n117), .Z(n115) );
  COND1XL U87 ( .A(n112), .B(n118), .C(n119), .Z(n648) );
  COND4CX1 U88 ( .A(\memory[27][2] ), .B(n45), .C(n120), .D(n112), .Z(n119) );
  COND2X1 U89 ( .A(n801), .B(n102), .C(n53), .D(n117), .Z(n120) );
  COND1XL U90 ( .A(n112), .B(n121), .C(n122), .Z(n649) );
  COND4CX1 U91 ( .A(\memory[27][1] ), .B(n45), .C(n123), .D(n112), .Z(n122) );
  COND2X1 U92 ( .A(n801), .B(n105), .C(n57), .D(n117), .Z(n123) );
  COND1XL U93 ( .A(n112), .B(n124), .C(n125), .Z(n650) );
  COND4CX1 U94 ( .A(\memory[27][0] ), .B(n45), .C(n126), .D(n112), .Z(n125) );
  COND2X1 U95 ( .A(n801), .B(n108), .C(n61), .D(n117), .Z(n126) );
  CANR1XL U96 ( .A(n117), .B(N282), .C(n62), .Z(n116) );
  COND1XL U97 ( .A(n39), .B(n117), .C(n16), .Z(n112) );
  CND2X1 U98 ( .A(n127), .B(n40), .Z(n117) );
  COND1XL U99 ( .A(n128), .B(n129), .C(n130), .Z(n651) );
  COND4CX1 U100 ( .A(\memory[26][3] ), .B(n45), .C(n131), .D(n128), .Z(n130)
         );
  COND2X1 U101 ( .A(n803), .B(n113), .C(n48), .D(n133), .Z(n131) );
  COND1XL U102 ( .A(n128), .B(n134), .C(n135), .Z(n652) );
  COND4CX1 U103 ( .A(\memory[26][2] ), .B(n45), .C(n136), .D(n128), .Z(n135)
         );
  COND2X1 U104 ( .A(n803), .B(n118), .C(n53), .D(n133), .Z(n136) );
  COND1XL U105 ( .A(n128), .B(n137), .C(n138), .Z(n653) );
  COND4CX1 U106 ( .A(\memory[26][1] ), .B(n45), .C(n139), .D(n128), .Z(n138)
         );
  COND2X1 U107 ( .A(n803), .B(n121), .C(n57), .D(n133), .Z(n139) );
  COND1XL U108 ( .A(n128), .B(n140), .C(n141), .Z(n654) );
  COND4CX1 U109 ( .A(\memory[26][0] ), .B(n45), .C(n142), .D(n128), .Z(n141)
         );
  COND2X1 U110 ( .A(n803), .B(n124), .C(n61), .D(n133), .Z(n142) );
  CANR1XL U111 ( .A(n133), .B(N282), .C(n62), .Z(n132) );
  COND1XL U112 ( .A(n39), .B(n133), .C(n16), .Z(n128) );
  CND2X1 U113 ( .A(n143), .B(n40), .Z(n133) );
  COND1XL U114 ( .A(n144), .B(n145), .C(n146), .Z(n655) );
  COND4CX1 U115 ( .A(\memory[25][3] ), .B(n45), .C(n147), .D(n144), .Z(n146)
         );
  COND2X1 U116 ( .A(n805), .B(n129), .C(n48), .D(n149), .Z(n147) );
  COND1XL U117 ( .A(n144), .B(n150), .C(n151), .Z(n656) );
  COND4CX1 U118 ( .A(\memory[25][2] ), .B(n45), .C(n152), .D(n144), .Z(n151)
         );
  COND2X1 U119 ( .A(n805), .B(n134), .C(n53), .D(n149), .Z(n152) );
  COND1XL U120 ( .A(n144), .B(n153), .C(n154), .Z(n657) );
  COND4CX1 U121 ( .A(\memory[25][1] ), .B(n45), .C(n155), .D(n144), .Z(n154)
         );
  COND2X1 U122 ( .A(n805), .B(n137), .C(n57), .D(n149), .Z(n155) );
  COND1XL U123 ( .A(n144), .B(n156), .C(n157), .Z(n658) );
  COND4CX1 U124 ( .A(\memory[25][0] ), .B(n45), .C(n158), .D(n144), .Z(n157)
         );
  COND2X1 U125 ( .A(n805), .B(n140), .C(n61), .D(n149), .Z(n158) );
  CANR1XL U126 ( .A(n149), .B(N282), .C(n62), .Z(n148) );
  COND1XL U127 ( .A(n39), .B(n149), .C(n16), .Z(n144) );
  CND2X1 U128 ( .A(n159), .B(n160), .Z(n149) );
  COND1XL U129 ( .A(n161), .B(n162), .C(n163), .Z(n659) );
  COND4CX1 U130 ( .A(\memory[24][3] ), .B(n45), .C(n164), .D(n161), .Z(n163)
         );
  COND2X1 U131 ( .A(n807), .B(n145), .C(n48), .D(n166), .Z(n164) );
  COND1XL U132 ( .A(n161), .B(n167), .C(n168), .Z(n660) );
  COND4CX1 U133 ( .A(\memory[24][2] ), .B(n45), .C(n169), .D(n161), .Z(n168)
         );
  COND2X1 U134 ( .A(n807), .B(n150), .C(n53), .D(n166), .Z(n169) );
  COND1XL U135 ( .A(n161), .B(n170), .C(n171), .Z(n661) );
  COND4CX1 U136 ( .A(\memory[24][1] ), .B(n45), .C(n172), .D(n161), .Z(n171)
         );
  COND2X1 U137 ( .A(n807), .B(n153), .C(n57), .D(n166), .Z(n172) );
  COND1XL U138 ( .A(n161), .B(n173), .C(n174), .Z(n662) );
  COND4CX1 U139 ( .A(\memory[24][0] ), .B(n45), .C(n175), .D(n161), .Z(n174)
         );
  COND2X1 U140 ( .A(n807), .B(n156), .C(n61), .D(n166), .Z(n175) );
  CANR1XL U141 ( .A(n166), .B(N282), .C(n62), .Z(n165) );
  COND1XL U142 ( .A(n39), .B(n166), .C(n16), .Z(n161) );
  CND2X1 U143 ( .A(n160), .B(n41), .Z(n166) );
  COND1XL U144 ( .A(n176), .B(n177), .C(n178), .Z(n663) );
  COND4CX1 U145 ( .A(\memory[23][3] ), .B(n45), .C(n179), .D(n176), .Z(n178)
         );
  COND2X1 U146 ( .A(n809), .B(n162), .C(n48), .D(n181), .Z(n179) );
  COND1XL U147 ( .A(n176), .B(n182), .C(n183), .Z(n664) );
  COND4CX1 U148 ( .A(\memory[23][2] ), .B(n45), .C(n184), .D(n176), .Z(n183)
         );
  COND2X1 U149 ( .A(n809), .B(n167), .C(n53), .D(n181), .Z(n184) );
  COND1XL U150 ( .A(n176), .B(n185), .C(n186), .Z(n665) );
  COND4CX1 U151 ( .A(\memory[23][1] ), .B(n45), .C(n187), .D(n176), .Z(n186)
         );
  COND2X1 U152 ( .A(n809), .B(n170), .C(n57), .D(n181), .Z(n187) );
  COND1XL U153 ( .A(n176), .B(n188), .C(n189), .Z(n666) );
  COND4CX1 U154 ( .A(\memory[23][0] ), .B(n45), .C(n190), .D(n176), .Z(n189)
         );
  COND2X1 U155 ( .A(n809), .B(n173), .C(n61), .D(n181), .Z(n190) );
  CANR1XL U156 ( .A(n181), .B(N282), .C(n62), .Z(n180) );
  COND1XL U157 ( .A(n39), .B(n181), .C(n16), .Z(n176) );
  CND2X1 U158 ( .A(n160), .B(n63), .Z(n181) );
  COND1XL U159 ( .A(n191), .B(n192), .C(n193), .Z(n667) );
  COND4CX1 U160 ( .A(\memory[22][3] ), .B(n45), .C(n194), .D(n191), .Z(n193)
         );
  COND2X1 U161 ( .A(n811), .B(n177), .C(n48), .D(n196), .Z(n194) );
  COND1XL U162 ( .A(n191), .B(n197), .C(n198), .Z(n668) );
  COND4CX1 U163 ( .A(\memory[22][2] ), .B(n45), .C(n199), .D(n191), .Z(n198)
         );
  COND2X1 U164 ( .A(n811), .B(n182), .C(n53), .D(n196), .Z(n199) );
  COND1XL U165 ( .A(n191), .B(n200), .C(n201), .Z(n669) );
  COND4CX1 U166 ( .A(\memory[22][1] ), .B(n45), .C(n202), .D(n191), .Z(n201)
         );
  COND2X1 U167 ( .A(n811), .B(n185), .C(n57), .D(n196), .Z(n202) );
  COND1XL U168 ( .A(n191), .B(n203), .C(n204), .Z(n670) );
  COND4CX1 U169 ( .A(\memory[22][0] ), .B(n45), .C(n205), .D(n191), .Z(n204)
         );
  COND2X1 U170 ( .A(n811), .B(n188), .C(n61), .D(n196), .Z(n205) );
  CANR1XL U171 ( .A(n196), .B(N282), .C(n62), .Z(n195) );
  COND1XL U172 ( .A(n39), .B(n196), .C(n16), .Z(n191) );
  CND2X1 U173 ( .A(n160), .B(n79), .Z(n196) );
  COND1XL U174 ( .A(n206), .B(n207), .C(n208), .Z(n671) );
  COND4CX1 U175 ( .A(\memory[21][3] ), .B(n45), .C(n209), .D(n206), .Z(n208)
         );
  COND2X1 U176 ( .A(n813), .B(n192), .C(n48), .D(n211), .Z(n209) );
  COND1XL U177 ( .A(n206), .B(n212), .C(n213), .Z(n672) );
  COND4CX1 U178 ( .A(\memory[21][2] ), .B(n45), .C(n214), .D(n206), .Z(n213)
         );
  COND2X1 U179 ( .A(n813), .B(n197), .C(n53), .D(n211), .Z(n214) );
  COND1XL U180 ( .A(n206), .B(n215), .C(n216), .Z(n673) );
  COND4CX1 U181 ( .A(\memory[21][1] ), .B(n45), .C(n217), .D(n206), .Z(n216)
         );
  COND2X1 U182 ( .A(n813), .B(n200), .C(n57), .D(n211), .Z(n217) );
  COND1XL U183 ( .A(n206), .B(n218), .C(n219), .Z(n674) );
  COND4CX1 U184 ( .A(\memory[21][0] ), .B(n45), .C(n220), .D(n206), .Z(n219)
         );
  COND2X1 U185 ( .A(n813), .B(n203), .C(n61), .D(n211), .Z(n220) );
  CANR1XL U186 ( .A(n211), .B(N282), .C(n62), .Z(n210) );
  COND1XL U187 ( .A(n39), .B(n211), .C(n16), .Z(n206) );
  CND2X1 U188 ( .A(n160), .B(n95), .Z(n211) );
  COND1XL U189 ( .A(n221), .B(n222), .C(n223), .Z(n675) );
  COND4CX1 U190 ( .A(\memory[20][3] ), .B(n45), .C(n224), .D(n221), .Z(n223)
         );
  COND2X1 U191 ( .A(n815), .B(n207), .C(n48), .D(n226), .Z(n224) );
  COND1XL U192 ( .A(n221), .B(n227), .C(n228), .Z(n676) );
  COND4CX1 U193 ( .A(\memory[20][2] ), .B(n45), .C(n229), .D(n221), .Z(n228)
         );
  COND2X1 U194 ( .A(n815), .B(n212), .C(n53), .D(n226), .Z(n229) );
  COND1XL U195 ( .A(n221), .B(n230), .C(n231), .Z(n677) );
  COND4CX1 U196 ( .A(\memory[20][1] ), .B(n45), .C(n232), .D(n221), .Z(n231)
         );
  COND2X1 U197 ( .A(n815), .B(n215), .C(n57), .D(n226), .Z(n232) );
  COND1XL U198 ( .A(n221), .B(n233), .C(n234), .Z(n678) );
  COND4CX1 U199 ( .A(\memory[20][0] ), .B(n45), .C(n235), .D(n221), .Z(n234)
         );
  COND2X1 U200 ( .A(n815), .B(n218), .C(n61), .D(n226), .Z(n235) );
  CANR1XL U201 ( .A(n226), .B(N282), .C(n62), .Z(n225) );
  COND1XL U202 ( .A(n39), .B(n226), .C(n16), .Z(n221) );
  CND2X1 U203 ( .A(n160), .B(n111), .Z(n226) );
  COND1XL U204 ( .A(n236), .B(n237), .C(n238), .Z(n679) );
  COND4CX1 U205 ( .A(\memory[19][3] ), .B(n45), .C(n239), .D(n236), .Z(n238)
         );
  COND2X1 U206 ( .A(n817), .B(n222), .C(n48), .D(n241), .Z(n239) );
  COND1XL U207 ( .A(n236), .B(n242), .C(n243), .Z(n680) );
  COND4CX1 U208 ( .A(\memory[19][2] ), .B(n45), .C(n244), .D(n236), .Z(n243)
         );
  COND2X1 U209 ( .A(n817), .B(n227), .C(n53), .D(n241), .Z(n244) );
  COND1XL U210 ( .A(n236), .B(n245), .C(n246), .Z(n681) );
  COND4CX1 U211 ( .A(\memory[19][1] ), .B(n45), .C(n247), .D(n236), .Z(n246)
         );
  COND2X1 U212 ( .A(n817), .B(n230), .C(n57), .D(n241), .Z(n247) );
  COND1XL U213 ( .A(n236), .B(n248), .C(n249), .Z(n682) );
  COND4CX1 U214 ( .A(\memory[19][0] ), .B(n45), .C(n250), .D(n236), .Z(n249)
         );
  COND2X1 U215 ( .A(n817), .B(n233), .C(n61), .D(n241), .Z(n250) );
  CANR1XL U216 ( .A(n241), .B(N282), .C(n62), .Z(n240) );
  COND1XL U217 ( .A(n39), .B(n241), .C(n16), .Z(n236) );
  CND2X1 U218 ( .A(n160), .B(n127), .Z(n241) );
  COND1XL U219 ( .A(n251), .B(n252), .C(n253), .Z(n683) );
  COND4CX1 U220 ( .A(\memory[18][3] ), .B(n45), .C(n254), .D(n251), .Z(n253)
         );
  COND2X1 U221 ( .A(n819), .B(n237), .C(n48), .D(n256), .Z(n254) );
  COND1XL U222 ( .A(n251), .B(n257), .C(n258), .Z(n684) );
  COND4CX1 U223 ( .A(\memory[18][2] ), .B(n45), .C(n259), .D(n251), .Z(n258)
         );
  COND2X1 U224 ( .A(n819), .B(n242), .C(n53), .D(n256), .Z(n259) );
  COND1XL U225 ( .A(n251), .B(n260), .C(n261), .Z(n685) );
  COND4CX1 U226 ( .A(\memory[18][1] ), .B(n45), .C(n262), .D(n251), .Z(n261)
         );
  COND2X1 U227 ( .A(n819), .B(n245), .C(n57), .D(n256), .Z(n262) );
  COND1XL U228 ( .A(n251), .B(n263), .C(n264), .Z(n686) );
  COND4CX1 U229 ( .A(\memory[18][0] ), .B(n45), .C(n265), .D(n251), .Z(n264)
         );
  COND2X1 U230 ( .A(n819), .B(n248), .C(n61), .D(n256), .Z(n265) );
  CANR1XL U231 ( .A(n256), .B(N282), .C(n62), .Z(n255) );
  COND1XL U232 ( .A(n39), .B(n256), .C(n16), .Z(n251) );
  CND2X1 U233 ( .A(n160), .B(n143), .Z(n256) );
  CNR2X1 U234 ( .A(n266), .B(N276), .Z(n160) );
  COND1XL U235 ( .A(n267), .B(n268), .C(n269), .Z(n687) );
  COND4CX1 U236 ( .A(\memory[17][3] ), .B(n45), .C(n270), .D(n267), .Z(n269)
         );
  COND2X1 U237 ( .A(n821), .B(n252), .C(n48), .D(n272), .Z(n270) );
  COND1XL U238 ( .A(n267), .B(n273), .C(n274), .Z(n688) );
  COND4CX1 U239 ( .A(\memory[17][2] ), .B(n45), .C(n275), .D(n267), .Z(n274)
         );
  COND2X1 U240 ( .A(n821), .B(n257), .C(n53), .D(n272), .Z(n275) );
  COND1XL U241 ( .A(n267), .B(n276), .C(n277), .Z(n689) );
  COND4CX1 U242 ( .A(\memory[17][1] ), .B(n45), .C(n278), .D(n267), .Z(n277)
         );
  COND2X1 U243 ( .A(n821), .B(n260), .C(n57), .D(n272), .Z(n278) );
  COND1XL U244 ( .A(n267), .B(n279), .C(n280), .Z(n690) );
  COND4CX1 U245 ( .A(\memory[17][0] ), .B(n45), .C(n281), .D(n267), .Z(n280)
         );
  COND2X1 U246 ( .A(n821), .B(n263), .C(n61), .D(n272), .Z(n281) );
  CANR1XL U247 ( .A(n272), .B(N282), .C(n62), .Z(n271) );
  COND1XL U248 ( .A(n39), .B(n272), .C(n16), .Z(n267) );
  CND2X1 U249 ( .A(n282), .B(n159), .Z(n272) );
  COND1XL U250 ( .A(n283), .B(n284), .C(n285), .Z(n691) );
  COND4CX1 U251 ( .A(\memory[16][3] ), .B(n45), .C(n286), .D(n283), .Z(n285)
         );
  COND2X1 U252 ( .A(n823), .B(n268), .C(n48), .D(n288), .Z(n286) );
  COND1XL U253 ( .A(n283), .B(n289), .C(n290), .Z(n692) );
  COND4CX1 U254 ( .A(\memory[16][2] ), .B(n45), .C(n291), .D(n283), .Z(n290)
         );
  COND2X1 U255 ( .A(n823), .B(n273), .C(n53), .D(n288), .Z(n291) );
  COND1XL U256 ( .A(n283), .B(n292), .C(n293), .Z(n693) );
  COND4CX1 U257 ( .A(\memory[16][1] ), .B(n45), .C(n294), .D(n283), .Z(n293)
         );
  COND2X1 U258 ( .A(n823), .B(n276), .C(n57), .D(n288), .Z(n294) );
  COND1XL U259 ( .A(n283), .B(n295), .C(n296), .Z(n694) );
  COND4CX1 U260 ( .A(\memory[16][0] ), .B(n45), .C(n297), .D(n283), .Z(n296)
         );
  COND2X1 U261 ( .A(n823), .B(n279), .C(n61), .D(n288), .Z(n297) );
  CANR1XL U262 ( .A(n288), .B(N282), .C(n62), .Z(n287) );
  COND1XL U263 ( .A(n39), .B(n288), .C(n16), .Z(n283) );
  CND2X1 U264 ( .A(n282), .B(n41), .Z(n288) );
  COND1XL U265 ( .A(n298), .B(n299), .C(n300), .Z(n695) );
  COND4CX1 U266 ( .A(\memory[15][3] ), .B(n45), .C(n301), .D(n298), .Z(n300)
         );
  COND2X1 U267 ( .A(n825), .B(n284), .C(n48), .D(n303), .Z(n301) );
  COND1XL U268 ( .A(n298), .B(n304), .C(n305), .Z(n696) );
  COND4CX1 U269 ( .A(\memory[15][2] ), .B(n45), .C(n306), .D(n298), .Z(n305)
         );
  COND2X1 U270 ( .A(n825), .B(n289), .C(n53), .D(n303), .Z(n306) );
  COND1XL U271 ( .A(n298), .B(n307), .C(n308), .Z(n697) );
  COND4CX1 U272 ( .A(\memory[15][1] ), .B(n45), .C(n309), .D(n298), .Z(n308)
         );
  COND2X1 U273 ( .A(n825), .B(n292), .C(n57), .D(n303), .Z(n309) );
  COND1XL U274 ( .A(n298), .B(n310), .C(n311), .Z(n698) );
  COND4CX1 U275 ( .A(\memory[15][0] ), .B(n45), .C(n312), .D(n298), .Z(n311)
         );
  COND2X1 U276 ( .A(n825), .B(n295), .C(n61), .D(n303), .Z(n312) );
  CANR1XL U277 ( .A(n303), .B(N282), .C(n62), .Z(n302) );
  COND1XL U278 ( .A(n39), .B(n303), .C(n16), .Z(n298) );
  CND2X1 U279 ( .A(n282), .B(n63), .Z(n303) );
  COND1XL U280 ( .A(n313), .B(n314), .C(n315), .Z(n699) );
  COND4CX1 U281 ( .A(\memory[14][3] ), .B(n45), .C(n316), .D(n313), .Z(n315)
         );
  COND2X1 U282 ( .A(n827), .B(n299), .C(n48), .D(n318), .Z(n316) );
  COND1XL U283 ( .A(n313), .B(n319), .C(n320), .Z(n700) );
  COND4CX1 U284 ( .A(\memory[14][2] ), .B(n45), .C(n321), .D(n313), .Z(n320)
         );
  COND2X1 U285 ( .A(n827), .B(n304), .C(n53), .D(n318), .Z(n321) );
  COND1XL U286 ( .A(n313), .B(n322), .C(n323), .Z(n701) );
  COND4CX1 U287 ( .A(\memory[14][1] ), .B(n45), .C(n324), .D(n313), .Z(n323)
         );
  COND2X1 U288 ( .A(n827), .B(n307), .C(n57), .D(n318), .Z(n324) );
  COND1XL U289 ( .A(n313), .B(n325), .C(n326), .Z(n702) );
  COND4CX1 U290 ( .A(\memory[14][0] ), .B(n45), .C(n327), .D(n313), .Z(n326)
         );
  COND2X1 U291 ( .A(n827), .B(n310), .C(n61), .D(n318), .Z(n327) );
  CANR1XL U292 ( .A(n318), .B(N282), .C(n62), .Z(n317) );
  COND1XL U293 ( .A(n39), .B(n318), .C(n16), .Z(n313) );
  CND2X1 U294 ( .A(n282), .B(n79), .Z(n318) );
  COND1XL U295 ( .A(n328), .B(n329), .C(n330), .Z(n703) );
  COND4CX1 U296 ( .A(\memory[13][3] ), .B(n45), .C(n331), .D(n328), .Z(n330)
         );
  COND2X1 U297 ( .A(n829), .B(n314), .C(n48), .D(n333), .Z(n331) );
  COND1XL U298 ( .A(n328), .B(n334), .C(n335), .Z(n704) );
  COND4CX1 U299 ( .A(\memory[13][2] ), .B(n45), .C(n336), .D(n328), .Z(n335)
         );
  COND2X1 U300 ( .A(n829), .B(n319), .C(n53), .D(n333), .Z(n336) );
  COND1XL U301 ( .A(n328), .B(n337), .C(n338), .Z(n705) );
  COND4CX1 U302 ( .A(\memory[13][1] ), .B(n45), .C(n339), .D(n328), .Z(n338)
         );
  COND2X1 U303 ( .A(n829), .B(n322), .C(n57), .D(n333), .Z(n339) );
  COND1XL U304 ( .A(n328), .B(n340), .C(n341), .Z(n706) );
  COND4CX1 U305 ( .A(\memory[13][0] ), .B(n45), .C(n342), .D(n328), .Z(n341)
         );
  COND2X1 U306 ( .A(n829), .B(n325), .C(n61), .D(n333), .Z(n342) );
  CANR1XL U307 ( .A(n333), .B(N282), .C(n62), .Z(n332) );
  COND1XL U308 ( .A(n39), .B(n333), .C(n16), .Z(n328) );
  CND2X1 U309 ( .A(n282), .B(n95), .Z(n333) );
  COND1XL U310 ( .A(n343), .B(n344), .C(n345), .Z(n707) );
  COND4CX1 U311 ( .A(\memory[12][3] ), .B(n45), .C(n346), .D(n343), .Z(n345)
         );
  COND2X1 U312 ( .A(n831), .B(n329), .C(n48), .D(n348), .Z(n346) );
  COND1XL U313 ( .A(n343), .B(n349), .C(n350), .Z(n708) );
  COND4CX1 U314 ( .A(\memory[12][2] ), .B(n45), .C(n351), .D(n343), .Z(n350)
         );
  COND2X1 U315 ( .A(n831), .B(n334), .C(n53), .D(n348), .Z(n351) );
  COND1XL U316 ( .A(n343), .B(n352), .C(n353), .Z(n709) );
  COND4CX1 U317 ( .A(\memory[12][1] ), .B(n45), .C(n354), .D(n343), .Z(n353)
         );
  COND2X1 U318 ( .A(n831), .B(n337), .C(n57), .D(n348), .Z(n354) );
  COND1XL U319 ( .A(n343), .B(n355), .C(n356), .Z(n710) );
  COND4CX1 U320 ( .A(\memory[12][0] ), .B(n45), .C(n357), .D(n343), .Z(n356)
         );
  COND2X1 U321 ( .A(n831), .B(n340), .C(n61), .D(n348), .Z(n357) );
  CANR1XL U322 ( .A(n348), .B(N282), .C(n62), .Z(n347) );
  COND1XL U323 ( .A(n39), .B(n348), .C(n16), .Z(n343) );
  CND2X1 U324 ( .A(n282), .B(n111), .Z(n348) );
  COND1XL U325 ( .A(n358), .B(n359), .C(n360), .Z(n711) );
  COND4CX1 U326 ( .A(\memory[11][3] ), .B(n45), .C(n361), .D(n358), .Z(n360)
         );
  COND2X1 U327 ( .A(n833), .B(n344), .C(n48), .D(n363), .Z(n361) );
  COND1XL U328 ( .A(n358), .B(n364), .C(n365), .Z(n712) );
  COND4CX1 U329 ( .A(\memory[11][2] ), .B(n45), .C(n366), .D(n358), .Z(n365)
         );
  COND2X1 U330 ( .A(n833), .B(n349), .C(n53), .D(n363), .Z(n366) );
  COND1XL U331 ( .A(n358), .B(n367), .C(n368), .Z(n713) );
  COND4CX1 U332 ( .A(\memory[11][1] ), .B(n45), .C(n369), .D(n358), .Z(n368)
         );
  COND2X1 U333 ( .A(n833), .B(n352), .C(n57), .D(n363), .Z(n369) );
  COND1XL U334 ( .A(n358), .B(n370), .C(n371), .Z(n714) );
  COND4CX1 U335 ( .A(\memory[11][0] ), .B(n45), .C(n372), .D(n358), .Z(n371)
         );
  COND2X1 U336 ( .A(n833), .B(n355), .C(n61), .D(n363), .Z(n372) );
  CANR1XL U337 ( .A(n363), .B(N282), .C(n62), .Z(n362) );
  COND1XL U338 ( .A(n39), .B(n363), .C(n16), .Z(n358) );
  CND2X1 U339 ( .A(n282), .B(n127), .Z(n363) );
  COND1XL U340 ( .A(n373), .B(n374), .C(n375), .Z(n715) );
  COND4CX1 U341 ( .A(\memory[10][3] ), .B(n45), .C(n376), .D(n373), .Z(n375)
         );
  COND2X1 U342 ( .A(n835), .B(n359), .C(n48), .D(n378), .Z(n376) );
  COND1XL U343 ( .A(n373), .B(n379), .C(n380), .Z(n716) );
  COND4CX1 U344 ( .A(\memory[10][2] ), .B(n45), .C(n381), .D(n373), .Z(n380)
         );
  COND2X1 U345 ( .A(n835), .B(n364), .C(n53), .D(n378), .Z(n381) );
  COND1XL U346 ( .A(n373), .B(n382), .C(n383), .Z(n717) );
  COND4CX1 U347 ( .A(\memory[10][1] ), .B(n45), .C(n384), .D(n373), .Z(n383)
         );
  COND2X1 U348 ( .A(n835), .B(n367), .C(n57), .D(n378), .Z(n384) );
  COND1XL U349 ( .A(n373), .B(n385), .C(n386), .Z(n718) );
  COND4CX1 U350 ( .A(\memory[10][0] ), .B(n45), .C(n387), .D(n373), .Z(n386)
         );
  COND2X1 U351 ( .A(n835), .B(n370), .C(n61), .D(n378), .Z(n387) );
  CANR1XL U352 ( .A(n378), .B(N282), .C(n62), .Z(n377) );
  COND1XL U353 ( .A(n39), .B(n378), .C(n16), .Z(n373) );
  CND2X1 U354 ( .A(n282), .B(n143), .Z(n378) );
  CNR2X1 U355 ( .A(n388), .B(N275), .Z(n282) );
  COND4CX1 U357 ( .A(\memory[9][3] ), .B(n45), .C(n392), .D(n389), .Z(n391) );
  COND2X1 U358 ( .A(n393), .B(n374), .C(n48), .D(n394), .Z(n392) );
  COND4CX1 U360 ( .A(\memory[9][2] ), .B(n45), .C(n397), .D(n389), .Z(n396) );
  COND2X1 U361 ( .A(n393), .B(n379), .C(n53), .D(n394), .Z(n397) );
  COND4CX1 U363 ( .A(\memory[9][1] ), .B(n45), .C(n400), .D(n389), .Z(n399) );
  COND2X1 U364 ( .A(n393), .B(n382), .C(n57), .D(n394), .Z(n400) );
  COND4CX1 U366 ( .A(\memory[9][0] ), .B(n45), .C(n403), .D(n389), .Z(n402) );
  COND2X1 U367 ( .A(n393), .B(n385), .C(n61), .D(n394), .Z(n403) );
  CANR1XL U368 ( .A(n394), .B(N282), .C(n62), .Z(n393) );
  COND1XL U369 ( .A(n39), .B(n394), .C(n16), .Z(n389) );
  CND2X1 U370 ( .A(n404), .B(n159), .Z(n394) );
  COND1XL U371 ( .A(n405), .B(n406), .C(n407), .Z(n723) );
  COND4CX1 U372 ( .A(\memory[8][3] ), .B(n45), .C(n408), .D(n405), .Z(n407) );
  COND2X1 U373 ( .A(n837), .B(n390), .C(n48), .D(n410), .Z(n408) );
  COND1XL U374 ( .A(n405), .B(n411), .C(n412), .Z(n724) );
  COND4CX1 U375 ( .A(\memory[8][2] ), .B(n45), .C(n413), .D(n405), .Z(n412) );
  COND2X1 U376 ( .A(n837), .B(n395), .C(n53), .D(n410), .Z(n413) );
  COND1XL U377 ( .A(n405), .B(n414), .C(n415), .Z(n725) );
  COND4CX1 U378 ( .A(\memory[8][1] ), .B(n45), .C(n416), .D(n405), .Z(n415) );
  COND2X1 U379 ( .A(n837), .B(n398), .C(n57), .D(n410), .Z(n416) );
  COND1XL U380 ( .A(n405), .B(n417), .C(n418), .Z(n726) );
  COND4CX1 U381 ( .A(\memory[8][0] ), .B(n45), .C(n419), .D(n405), .Z(n418) );
  COND2X1 U382 ( .A(n837), .B(n401), .C(n61), .D(n410), .Z(n419) );
  CANR1XL U383 ( .A(n410), .B(N282), .C(n62), .Z(n409) );
  COND1XL U384 ( .A(n39), .B(n410), .C(n16), .Z(n405) );
  CND2X1 U385 ( .A(n404), .B(n41), .Z(n410) );
  CNR3XL U386 ( .A(n420), .B(N279), .C(n421), .Z(n41) );
  COND4CX1 U388 ( .A(\memory[7][3] ), .B(n45), .C(n425), .D(n422), .Z(n424) );
  COND2X1 U389 ( .A(n426), .B(n406), .C(n48), .D(n427), .Z(n425) );
  COND4CX1 U391 ( .A(\memory[7][2] ), .B(n45), .C(n430), .D(n422), .Z(n429) );
  COND2X1 U392 ( .A(n426), .B(n411), .C(n53), .D(n427), .Z(n430) );
  COND4CX1 U394 ( .A(\memory[7][1] ), .B(n45), .C(n433), .D(n422), .Z(n432) );
  COND2X1 U395 ( .A(n426), .B(n414), .C(n57), .D(n427), .Z(n433) );
  COND4CX1 U397 ( .A(\memory[7][0] ), .B(n45), .C(n436), .D(n422), .Z(n435) );
  COND2X1 U398 ( .A(n426), .B(n417), .C(n61), .D(n427), .Z(n436) );
  CANR1XL U399 ( .A(n427), .B(N282), .C(n62), .Z(n426) );
  COND1XL U400 ( .A(n39), .B(n427), .C(n16), .Z(n422) );
  CND2X1 U401 ( .A(n404), .B(n63), .Z(n427) );
  CNR3XL U402 ( .A(n437), .B(N278), .C(n421), .Z(n63) );
  COND4CX1 U404 ( .A(\memory[6][3] ), .B(n45), .C(n441), .D(n438), .Z(n440) );
  COND2X1 U405 ( .A(n442), .B(n423), .C(n48), .D(n443), .Z(n441) );
  COND4CX1 U407 ( .A(\memory[6][2] ), .B(n45), .C(n446), .D(n438), .Z(n445) );
  COND2X1 U408 ( .A(n442), .B(n428), .C(n53), .D(n443), .Z(n446) );
  COND4CX1 U410 ( .A(\memory[6][1] ), .B(n45), .C(n449), .D(n438), .Z(n448) );
  COND2X1 U411 ( .A(n442), .B(n431), .C(n57), .D(n443), .Z(n449) );
  COND4CX1 U413 ( .A(\memory[6][0] ), .B(n45), .C(n452), .D(n438), .Z(n451) );
  COND2X1 U414 ( .A(n442), .B(n434), .C(n61), .D(n443), .Z(n452) );
  CANR1XL U415 ( .A(n443), .B(N282), .C(n62), .Z(n442) );
  COND1XL U416 ( .A(n39), .B(n443), .C(n16), .Z(n438) );
  CND2X1 U417 ( .A(n404), .B(n79), .Z(n443) );
  CNR3XL U418 ( .A(N278), .B(N279), .C(n421), .Z(n79) );
  COND4CX1 U420 ( .A(\memory[5][3] ), .B(n45), .C(n456), .D(n453), .Z(n455) );
  COND2X1 U421 ( .A(n457), .B(n439), .C(n48), .D(n458), .Z(n456) );
  COND4CX1 U423 ( .A(\memory[5][2] ), .B(n45), .C(n461), .D(n453), .Z(n460) );
  COND2X1 U424 ( .A(n457), .B(n444), .C(n53), .D(n458), .Z(n461) );
  COND4CX1 U426 ( .A(\memory[5][1] ), .B(n45), .C(n464), .D(n453), .Z(n463) );
  COND2X1 U427 ( .A(n457), .B(n447), .C(n57), .D(n458), .Z(n464) );
  COND4CX1 U429 ( .A(\memory[5][0] ), .B(n45), .C(n467), .D(n453), .Z(n466) );
  COND2X1 U430 ( .A(n457), .B(n450), .C(n61), .D(n458), .Z(n467) );
  CANR1XL U431 ( .A(n458), .B(N282), .C(n62), .Z(n457) );
  COND1XL U432 ( .A(n39), .B(n458), .C(n16), .Z(n453) );
  CND2X1 U433 ( .A(n404), .B(n95), .Z(n458) );
  CNR3XL U434 ( .A(n437), .B(N277), .C(n420), .Z(n95) );
  COND4CX1 U436 ( .A(\memory[4][3] ), .B(n45), .C(n471), .D(n468), .Z(n470) );
  COND2X1 U437 ( .A(n472), .B(n454), .C(n48), .D(n473), .Z(n471) );
  COND4CX1 U439 ( .A(\memory[4][2] ), .B(n45), .C(n476), .D(n468), .Z(n475) );
  COND2X1 U440 ( .A(n472), .B(n459), .C(n53), .D(n473), .Z(n476) );
  COND4CX1 U442 ( .A(\memory[4][1] ), .B(n45), .C(n479), .D(n468), .Z(n478) );
  COND2X1 U443 ( .A(n472), .B(n462), .C(n57), .D(n473), .Z(n479) );
  COND4CX1 U445 ( .A(\memory[4][0] ), .B(n45), .C(n482), .D(n468), .Z(n481) );
  COND2X1 U446 ( .A(n472), .B(n465), .C(n61), .D(n473), .Z(n482) );
  CANR1XL U447 ( .A(n473), .B(N282), .C(n62), .Z(n472) );
  COND1XL U448 ( .A(n39), .B(n473), .C(n16), .Z(n468) );
  CND2X1 U449 ( .A(n404), .B(n111), .Z(n473) );
  CNR3XL U450 ( .A(N277), .B(N279), .C(n420), .Z(n111) );
  COND4CX1 U452 ( .A(\memory[3][3] ), .B(n45), .C(n486), .D(n483), .Z(n485) );
  COND2X1 U453 ( .A(n487), .B(n469), .C(n48), .D(n488), .Z(n486) );
  COND4CX1 U455 ( .A(\memory[3][2] ), .B(n45), .C(n491), .D(n483), .Z(n490) );
  COND2X1 U456 ( .A(n487), .B(n474), .C(n53), .D(n488), .Z(n491) );
  COND4CX1 U458 ( .A(\memory[3][1] ), .B(n45), .C(n494), .D(n483), .Z(n493) );
  COND2X1 U459 ( .A(n487), .B(n477), .C(n57), .D(n488), .Z(n494) );
  COND2X1 U462 ( .A(n487), .B(n480), .C(n61), .D(n488), .Z(n497) );
  CANR1XL U463 ( .A(n488), .B(N282), .C(n62), .Z(n487) );
  COND1XL U464 ( .A(n39), .B(n488), .C(n16), .Z(n483) );
  CND2X1 U465 ( .A(n404), .B(n127), .Z(n488) );
  CNR3XL U466 ( .A(N277), .B(N278), .C(n437), .Z(n127) );
  CAOR2X1 U467 ( .A(code[3]), .B(n498), .C(\memory[0][3] ), .D(n499), .Z(n747)
         );
  COND1XL U468 ( .A(n500), .B(n501), .C(n502), .Z(n748) );
  COND4CX1 U469 ( .A(\memory[2][3] ), .B(n45), .C(n503), .D(n501), .Z(n502) );
  COND2X1 U470 ( .A(n791), .B(n484), .C(n48), .D(n505), .Z(n503) );
  CIVX1 U471 ( .A(n27), .Z(n48) );
  CNR2IX1 U472 ( .B(data[3]), .A(n21), .Z(n27) );
  CAOR2X1 U474 ( .A(code[2]), .B(n498), .C(\memory[0][2] ), .D(n499), .Z(n749)
         );
  COND1XL U475 ( .A(n501), .B(n506), .C(n507), .Z(n750) );
  COND4CX1 U476 ( .A(\memory[2][2] ), .B(n45), .C(n508), .D(n501), .Z(n507) );
  COND2X1 U477 ( .A(n791), .B(n489), .C(n53), .D(n505), .Z(n508) );
  CIVX1 U478 ( .A(n31), .Z(n53) );
  CNR2IX1 U479 ( .B(data[2]), .A(n21), .Z(n31) );
  CAOR2X1 U481 ( .A(code[1]), .B(n498), .C(\memory[0][1] ), .D(n499), .Z(n751)
         );
  COND1XL U482 ( .A(n501), .B(n509), .C(n510), .Z(n752) );
  COND4CX1 U483 ( .A(\memory[2][1] ), .B(n45), .C(n511), .D(n501), .Z(n510) );
  COND2X1 U484 ( .A(n791), .B(n492), .C(n57), .D(n505), .Z(n511) );
  CIVX1 U485 ( .A(n34), .Z(n57) );
  CNR2IX1 U486 ( .B(data[1]), .A(n21), .Z(n34) );
  CAOR2X1 U488 ( .A(code[0]), .B(n498), .C(\memory[0][0] ), .D(n499), .Z(n753)
         );
  CIVX1 U489 ( .A(n498), .Z(n499) );
  COND1XL U490 ( .A(n501), .B(n512), .C(n513), .Z(n754) );
  COND4CX1 U491 ( .A(\memory[2][0] ), .B(n45), .C(n514), .D(n501), .Z(n513) );
  COND2X1 U492 ( .A(n791), .B(n495), .C(n61), .D(n505), .Z(n514) );
  CIVX1 U493 ( .A(n37), .Z(n61) );
  CNR2IX1 U494 ( .B(data[0]), .A(n21), .Z(n37) );
  CANR1XL U495 ( .A(n505), .B(N282), .C(n62), .Z(n504) );
  COND1XL U496 ( .A(N282), .B(n515), .C(wr_enable), .Z(n62) );
  COND1XL U499 ( .A(n39), .B(n505), .C(n16), .Z(n501) );
  CIVX1 U500 ( .A(n18), .Z(n16) );
  COND1XL U501 ( .A(N282), .B(n39), .C(n498), .Z(n18) );
  CNR3XL U503 ( .A(n516), .B(n517), .C(n518), .Z(n515) );
  CND2X1 U505 ( .A(n404), .B(n143), .Z(n505) );
  CNR3XL U506 ( .A(N278), .B(N279), .C(N277), .Z(n143) );
  CNR2X1 U507 ( .A(N275), .B(N276), .Z(n404) );
  CAOR2X1 U508 ( .A(data[3]), .B(n519), .C(n520), .D(\memory[31][3] ), .Z(n755) );
  CAOR2X1 U509 ( .A(data[2]), .B(n519), .C(n520), .D(\memory[31][2] ), .Z(n756) );
  CAOR2X1 U510 ( .A(data[1]), .B(n519), .C(n520), .D(\memory[31][1] ), .Z(n757) );
  CAOR2X1 U511 ( .A(data[0]), .B(n519), .C(n520), .D(\memory[31][0] ), .Z(n758) );
  CIVX1 U512 ( .A(n520), .Z(n519) );
  COND4CX1 U513 ( .A(n159), .B(n40), .C(n521), .D(n522), .Z(n520) );
  CIVX1 U514 ( .A(n39), .Z(n522) );
  CND2X1 U515 ( .A(wr_enable), .B(reset), .Z(n39) );
  CNR2X1 U517 ( .A(n266), .B(n388), .Z(n40) );
  CNR3XL U518 ( .A(n420), .B(n437), .C(n421), .Z(n159) );
  CND2X1 U521 ( .A(N593), .B(n529), .Z(n525) );
  COND3X1 U522 ( .A(n530), .B(n524), .C(n531), .D(n532), .Z(n760) );
  CANR2X1 U523 ( .A(N119), .B(n527), .C(counter[29]), .D(n528), .Z(n532) );
  CND2X1 U524 ( .A(N592), .B(n529), .Z(n531) );
  CANR2X1 U526 ( .A(N117), .B(n527), .C(counter[28]), .D(n528), .Z(n535) );
  CND2X1 U527 ( .A(N591), .B(n529), .Z(n534) );
  COND3X1 U528 ( .A(n536), .B(n524), .C(n537), .D(n538), .Z(n762) );
  CANR2X1 U529 ( .A(N115), .B(n527), .C(counter[27]), .D(n528), .Z(n538) );
  CND2X1 U530 ( .A(N590), .B(n529), .Z(n537) );
  COND3X1 U531 ( .A(n539), .B(n524), .C(n540), .D(n541), .Z(n763) );
  CANR2X1 U532 ( .A(N113), .B(n527), .C(counter[26]), .D(n528), .Z(n541) );
  CND2X1 U533 ( .A(N589), .B(n529), .Z(n540) );
  COND3X1 U534 ( .A(n542), .B(n524), .C(n543), .D(n544), .Z(n764) );
  CANR2X1 U535 ( .A(N111), .B(n527), .C(counter[25]), .D(n528), .Z(n544) );
  CND2X1 U536 ( .A(N588), .B(n529), .Z(n543) );
  COND3X1 U537 ( .A(n545), .B(n524), .C(n546), .D(n547), .Z(n765) );
  CANR2X1 U538 ( .A(N109), .B(n527), .C(counter[24]), .D(n528), .Z(n547) );
  CND2X1 U539 ( .A(N587), .B(n529), .Z(n546) );
  COND3X1 U540 ( .A(n548), .B(n524), .C(n549), .D(n550), .Z(n766) );
  CANR2X1 U541 ( .A(N107), .B(n527), .C(counter[23]), .D(n528), .Z(n550) );
  CND2X1 U542 ( .A(N586), .B(n529), .Z(n549) );
  COND3X1 U543 ( .A(n551), .B(n524), .C(n552), .D(n553), .Z(n767) );
  CANR2X1 U544 ( .A(N105), .B(n527), .C(counter[22]), .D(n528), .Z(n553) );
  CND2X1 U545 ( .A(N585), .B(n529), .Z(n552) );
  COND3X1 U546 ( .A(n554), .B(n524), .C(n555), .D(n556), .Z(n768) );
  CANR2X1 U547 ( .A(N103), .B(n527), .C(counter[21]), .D(n528), .Z(n556) );
  CND2X1 U548 ( .A(N584), .B(n529), .Z(n555) );
  COND3X1 U549 ( .A(n557), .B(n524), .C(n558), .D(n559), .Z(n769) );
  CANR2X1 U550 ( .A(N101), .B(n527), .C(counter[20]), .D(n528), .Z(n559) );
  CND2X1 U551 ( .A(N583), .B(n529), .Z(n558) );
  COND3X1 U552 ( .A(n560), .B(n524), .C(n561), .D(n562), .Z(n770) );
  CANR2X1 U553 ( .A(N99), .B(n527), .C(counter[19]), .D(n528), .Z(n562) );
  CND2X1 U554 ( .A(N582), .B(n529), .Z(n561) );
  COND3X1 U555 ( .A(n563), .B(n524), .C(n564), .D(n565), .Z(n771) );
  CANR2X1 U556 ( .A(N97), .B(n527), .C(counter[18]), .D(n528), .Z(n565) );
  CND2X1 U557 ( .A(N581), .B(n529), .Z(n564) );
  COND3X1 U558 ( .A(n566), .B(n524), .C(n567), .D(n568), .Z(n772) );
  CANR2X1 U559 ( .A(N95), .B(n527), .C(counter[17]), .D(n528), .Z(n568) );
  CND2X1 U560 ( .A(N580), .B(n529), .Z(n567) );
  COND3X1 U561 ( .A(n569), .B(n524), .C(n570), .D(n571), .Z(n773) );
  CANR2X1 U562 ( .A(N93), .B(n527), .C(counter[16]), .D(n528), .Z(n571) );
  CND2X1 U563 ( .A(N579), .B(n529), .Z(n570) );
  COND3X1 U564 ( .A(n572), .B(n524), .C(n573), .D(n574), .Z(n774) );
  CANR2X1 U565 ( .A(N91), .B(n527), .C(counter[15]), .D(n528), .Z(n574) );
  CND2X1 U566 ( .A(N578), .B(n529), .Z(n573) );
  COND3X1 U567 ( .A(n575), .B(n524), .C(n576), .D(n577), .Z(n775) );
  CANR2X1 U568 ( .A(N89), .B(n527), .C(counter[14]), .D(n528), .Z(n577) );
  CND2X1 U569 ( .A(N577), .B(n529), .Z(n576) );
  COND3X1 U570 ( .A(n578), .B(n524), .C(n579), .D(n580), .Z(n776) );
  CANR2X1 U571 ( .A(N87), .B(n527), .C(counter[13]), .D(n528), .Z(n580) );
  CND2X1 U572 ( .A(N576), .B(n529), .Z(n579) );
  COND3X1 U573 ( .A(n581), .B(n524), .C(n582), .D(n583), .Z(n777) );
  CANR2X1 U574 ( .A(N85), .B(n527), .C(counter[12]), .D(n528), .Z(n583) );
  CND2X1 U575 ( .A(N575), .B(n529), .Z(n582) );
  COND3X1 U576 ( .A(n584), .B(n524), .C(n585), .D(n586), .Z(n778) );
  CANR2X1 U577 ( .A(N83), .B(n527), .C(counter[11]), .D(n528), .Z(n586) );
  CND2X1 U578 ( .A(N574), .B(n529), .Z(n585) );
  COND3X1 U579 ( .A(n587), .B(n524), .C(n588), .D(n589), .Z(n779) );
  CANR2X1 U580 ( .A(N81), .B(n527), .C(counter[10]), .D(n528), .Z(n589) );
  CND2X1 U581 ( .A(N573), .B(n529), .Z(n588) );
  COND3X1 U582 ( .A(n590), .B(n524), .C(n591), .D(n592), .Z(n780) );
  CANR2X1 U583 ( .A(N79), .B(n527), .C(counter[9]), .D(n528), .Z(n592) );
  CND2X1 U584 ( .A(N572), .B(n529), .Z(n591) );
  COND3X1 U585 ( .A(n593), .B(n524), .C(n594), .D(n595), .Z(n781) );
  CANR2X1 U586 ( .A(N77), .B(n527), .C(counter[8]), .D(n528), .Z(n595) );
  CND2X1 U587 ( .A(N571), .B(n529), .Z(n594) );
  COND3X1 U588 ( .A(n596), .B(n524), .C(n597), .D(n598), .Z(n782) );
  CANR2X1 U589 ( .A(N75), .B(n527), .C(counter[7]), .D(n528), .Z(n598) );
  CND2X1 U590 ( .A(N570), .B(n529), .Z(n597) );
  COND3X1 U591 ( .A(n599), .B(n524), .C(n600), .D(n601), .Z(n783) );
  CANR2X1 U592 ( .A(N73), .B(n527), .C(counter[6]), .D(n528), .Z(n601) );
  CND2X1 U593 ( .A(N569), .B(n529), .Z(n600) );
  COND3X1 U594 ( .A(n602), .B(n524), .C(n603), .D(n604), .Z(n784) );
  CANR2X1 U595 ( .A(N71), .B(n527), .C(counter[5]), .D(n528), .Z(n604) );
  CND2X1 U596 ( .A(N568), .B(n529), .Z(n603) );
  COND3X1 U597 ( .A(n266), .B(n524), .C(n605), .D(n606), .Z(n785) );
  CANR2X1 U598 ( .A(n527), .B(N69), .C(counter[4]), .D(n528), .Z(n606) );
  CND2X1 U599 ( .A(N567), .B(n529), .Z(n605) );
  COND3X1 U600 ( .A(n388), .B(n524), .C(n607), .D(n608), .Z(n786) );
  CANR2X1 U601 ( .A(n527), .B(N67), .C(counter[3]), .D(n528), .Z(n608) );
  CND2X1 U602 ( .A(N566), .B(n529), .Z(n607) );
  COND3X1 U603 ( .A(n421), .B(n524), .C(n609), .D(n610), .Z(n787) );
  CANR2X1 U604 ( .A(n527), .B(N65), .C(counter[2]), .D(n528), .Z(n610) );
  CND2X1 U605 ( .A(N565), .B(n529), .Z(n609) );
  COND3X1 U606 ( .A(n420), .B(n524), .C(n611), .D(n612), .Z(n788) );
  CANR2X1 U607 ( .A(n527), .B(N63), .C(counter[1]), .D(n528), .Z(n612) );
  CND2X1 U608 ( .A(N564), .B(n529), .Z(n611) );
  CND2X1 U611 ( .A(N594), .B(n529), .Z(n614) );
  COND3X1 U612 ( .A(n437), .B(n524), .C(n616), .D(n617), .Z(n790) );
  CANR2X1 U613 ( .A(n527), .B(N61), .C(n14), .D(n528), .Z(n617) );
  CND2X1 U615 ( .A(N563), .B(n529), .Z(n616) );
  CND2X1 U617 ( .A(N282), .B(wr_enable), .Z(n21) );
  CND2X1 U619 ( .A(n618), .B(n619), .Z(n524) );
  CIVX1 U622 ( .A(wr_enable), .Z(n619) );
  CIVX1 U623 ( .A(n437), .Z(N279) );
  CANR2X1 U624 ( .A(n22), .B(N61), .C(n620), .D(n14), .Z(n437) );
  CIVX1 U625 ( .A(n420), .Z(N278) );
  CANR2X1 U626 ( .A(n22), .B(N63), .C(n620), .D(counter[1]), .Z(n420) );
  CIVX1 U627 ( .A(n421), .Z(N277) );
  CANR2X1 U628 ( .A(n22), .B(N65), .C(n620), .D(counter[2]), .Z(n421) );
  CIVX1 U629 ( .A(n388), .Z(N276) );
  CANR2X1 U630 ( .A(n22), .B(N67), .C(n620), .D(counter[3]), .Z(n388) );
  CIVX1 U631 ( .A(n266), .Z(N275) );
  CANR2X1 U632 ( .A(n22), .B(N69), .C(n620), .D(counter[4]), .Z(n266) );
  CIVX1 U633 ( .A(n602), .Z(N274) );
  CANR2X1 U634 ( .A(n22), .B(N71), .C(n620), .D(counter[5]), .Z(n602) );
  CIVX1 U635 ( .A(n599), .Z(N273) );
  CANR2X1 U636 ( .A(n22), .B(N73), .C(n620), .D(counter[6]), .Z(n599) );
  CIVX1 U637 ( .A(n596), .Z(N272) );
  CANR2X1 U638 ( .A(n22), .B(N75), .C(n620), .D(counter[7]), .Z(n596) );
  CIVX1 U639 ( .A(n593), .Z(N271) );
  CANR2X1 U640 ( .A(n22), .B(N77), .C(n620), .D(counter[8]), .Z(n593) );
  CIVX1 U641 ( .A(n590), .Z(N270) );
  CANR2X1 U642 ( .A(n22), .B(N79), .C(n620), .D(counter[9]), .Z(n590) );
  CIVX1 U643 ( .A(n587), .Z(N269) );
  CANR2X1 U644 ( .A(n22), .B(N81), .C(n620), .D(counter[10]), .Z(n587) );
  CIVX1 U645 ( .A(n584), .Z(N268) );
  CANR2X1 U646 ( .A(n22), .B(N83), .C(n620), .D(counter[11]), .Z(n584) );
  CIVX1 U647 ( .A(n581), .Z(N267) );
  CANR2X1 U648 ( .A(n22), .B(N85), .C(n620), .D(counter[12]), .Z(n581) );
  CIVX1 U649 ( .A(n578), .Z(N266) );
  CANR2X1 U650 ( .A(n22), .B(N87), .C(n620), .D(counter[13]), .Z(n578) );
  CIVX1 U651 ( .A(n575), .Z(N265) );
  CANR2X1 U652 ( .A(n22), .B(N89), .C(n620), .D(counter[14]), .Z(n575) );
  CIVX1 U653 ( .A(n572), .Z(N264) );
  CANR2X1 U654 ( .A(n22), .B(N91), .C(n620), .D(counter[15]), .Z(n572) );
  CIVX1 U655 ( .A(n569), .Z(N263) );
  CANR2X1 U656 ( .A(n22), .B(N93), .C(n620), .D(counter[16]), .Z(n569) );
  CIVX1 U657 ( .A(n566), .Z(N262) );
  CANR2X1 U658 ( .A(n22), .B(N95), .C(n620), .D(counter[17]), .Z(n566) );
  CIVX1 U659 ( .A(n563), .Z(N261) );
  CANR2X1 U660 ( .A(n22), .B(N97), .C(n620), .D(counter[18]), .Z(n563) );
  CIVX1 U661 ( .A(n560), .Z(N260) );
  CANR2X1 U662 ( .A(n22), .B(N99), .C(n620), .D(counter[19]), .Z(n560) );
  CIVX1 U663 ( .A(n557), .Z(N259) );
  CANR2X1 U664 ( .A(n22), .B(N101), .C(n620), .D(counter[20]), .Z(n557) );
  CIVX1 U665 ( .A(n554), .Z(N258) );
  CANR2X1 U666 ( .A(n22), .B(N103), .C(n620), .D(counter[21]), .Z(n554) );
  CIVX1 U667 ( .A(n551), .Z(N257) );
  CANR2X1 U668 ( .A(n22), .B(N105), .C(n620), .D(counter[22]), .Z(n551) );
  CIVX1 U669 ( .A(n548), .Z(N256) );
  CANR2X1 U670 ( .A(n22), .B(N107), .C(n620), .D(counter[23]), .Z(n548) );
  CIVX1 U671 ( .A(n545), .Z(N255) );
  CANR2X1 U672 ( .A(n22), .B(N109), .C(n620), .D(counter[24]), .Z(n545) );
  CIVX1 U673 ( .A(n542), .Z(N254) );
  CANR2X1 U674 ( .A(n22), .B(N111), .C(n620), .D(counter[25]), .Z(n542) );
  CIVX1 U675 ( .A(n539), .Z(N253) );
  CANR2X1 U676 ( .A(n22), .B(N113), .C(n620), .D(counter[26]), .Z(n539) );
  CIVX1 U677 ( .A(n536), .Z(N252) );
  CANR2X1 U678 ( .A(n22), .B(N115), .C(n620), .D(counter[27]), .Z(n536) );
  CIVX1 U679 ( .A(n533), .Z(N251) );
  CANR2X1 U680 ( .A(n22), .B(N117), .C(n620), .D(counter[28]), .Z(n533) );
  CIVX1 U681 ( .A(n530), .Z(N250) );
  CANR2X1 U682 ( .A(n22), .B(N119), .C(n620), .D(counter[29]), .Z(n530) );
  CIVX1 U683 ( .A(n523), .Z(N249) );
  CANR2X1 U684 ( .A(N121), .B(n22), .C(n620), .D(counter[30]), .Z(n523) );
  CIVX1 U687 ( .A(n22), .Z(n620) );
  CIVX1 U689 ( .A(N50), .Z(n516) );
  CAN4X1 U690 ( .A(n621), .B(n622), .C(n623), .D(n624), .Z(n517) );
  CNR8X1 U691 ( .A(counter[31]), .B(counter[3]), .C(counter[4]), .D(counter[5]), .E(counter[6]), .F(counter[7]), .G(counter[8]), .H(counter[9]), .Z(n624) );
  CNR8X1 U692 ( .A(counter[24]), .B(counter[25]), .C(counter[26]), .D(
        counter[27]), .E(counter[28]), .F(counter[29]), .G(counter[2]), .H(
        counter[30]), .Z(n623) );
  CNR8X1 U693 ( .A(counter[17]), .B(counter[18]), .C(counter[19]), .D(
        counter[1]), .E(counter[20]), .F(counter[21]), .G(counter[22]), .H(
        counter[23]), .Z(n622) );
  CNR8X1 U694 ( .A(n14), .B(counter[10]), .C(counter[11]), .D(counter[12]), 
        .E(counter[13]), .F(counter[14]), .G(counter[15]), .H(counter[16]), 
        .Z(n621) );
  CIVX1 U695 ( .A(reset), .Z(N1652) );
  CFD1XL \memory_reg[0][3]  ( .D(n748), .CP(clock), .Q(\memory[0][3] ), .QN(
        n500) );
  CFD1XL \memory_reg[0][2]  ( .D(n750), .CP(clock), .Q(\memory[0][2] ), .QN(
        n506) );
  CFD1XL \memory_reg[0][1]  ( .D(n752), .CP(clock), .Q(\memory[0][1] ), .QN(
        n509) );
  CFD1XL \memory_reg[0][0]  ( .D(n754), .CP(clock), .Q(\memory[0][0] ), .QN(
        n512) );
  CFD1XL \memory_reg[1][3]  ( .D(n743), .CP(clock), .QN(n484) );
  CFD1XL \memory_reg[1][2]  ( .D(n744), .CP(clock), .QN(n489) );
  CFD1XL \memory_reg[1][1]  ( .D(n745), .CP(clock), .QN(n492) );
  CFD1XL \memory_reg[1][0]  ( .D(n746), .CP(clock), .QN(n495) );
  CFD1XL \memory_reg[30][3]  ( .D(n627), .CP(clock), .Q(\memory[30][3] ), .QN(
        n24) );
  CFD1XL \memory_reg[30][2]  ( .D(n628), .CP(clock), .Q(\memory[30][2] ), .QN(
        n29) );
  CFD1XL \memory_reg[30][1]  ( .D(n629), .CP(clock), .Q(\memory[30][1] ), .QN(
        n32) );
  CFD1XL \memory_reg[30][0]  ( .D(n630), .CP(clock), .Q(\memory[30][0] ), .QN(
        n35) );
  CFD1XL \memory_reg[29][3]  ( .D(n631), .CP(clock), .Q(\memory[29][3] ), .QN(
        n43) );
  CFD1XL \memory_reg[29][2]  ( .D(n632), .CP(clock), .Q(\memory[29][2] ), .QN(
        n50) );
  CFD1XL \memory_reg[29][1]  ( .D(n633), .CP(clock), .Q(\memory[29][1] ), .QN(
        n54) );
  CFD1XL \memory_reg[29][0]  ( .D(n634), .CP(clock), .Q(\memory[29][0] ), .QN(
        n58) );
  CFD1XL \memory_reg[28][3]  ( .D(n635), .CP(clock), .Q(\memory[28][3] ), .QN(
        n65) );
  CFD1XL \memory_reg[28][2]  ( .D(n636), .CP(clock), .Q(\memory[28][2] ), .QN(
        n70) );
  CFD1XL \memory_reg[28][1]  ( .D(n637), .CP(clock), .Q(\memory[28][1] ), .QN(
        n73) );
  CFD1XL \memory_reg[28][0]  ( .D(n638), .CP(clock), .Q(\memory[28][0] ), .QN(
        n76) );
  CFD1XL \memory_reg[27][3]  ( .D(n639), .CP(clock), .Q(\memory[27][3] ), .QN(
        n81) );
  CFD1XL \memory_reg[27][2]  ( .D(n640), .CP(clock), .Q(\memory[27][2] ), .QN(
        n86) );
  CFD1XL \memory_reg[27][1]  ( .D(n641), .CP(clock), .Q(\memory[27][1] ), .QN(
        n89) );
  CFD1XL \memory_reg[27][0]  ( .D(n642), .CP(clock), .Q(\memory[27][0] ), .QN(
        n92) );
  CFD1XL \memory_reg[26][3]  ( .D(n643), .CP(clock), .Q(\memory[26][3] ), .QN(
        n97) );
  CFD1XL \memory_reg[26][2]  ( .D(n644), .CP(clock), .Q(\memory[26][2] ), .QN(
        n102) );
  CFD1XL \memory_reg[26][1]  ( .D(n645), .CP(clock), .Q(\memory[26][1] ), .QN(
        n105) );
  CFD1XL \memory_reg[26][0]  ( .D(n646), .CP(clock), .Q(\memory[26][0] ), .QN(
        n108) );
  CFD1XL \memory_reg[25][3]  ( .D(n647), .CP(clock), .Q(\memory[25][3] ), .QN(
        n113) );
  CFD1XL \memory_reg[25][2]  ( .D(n648), .CP(clock), .Q(\memory[25][2] ), .QN(
        n118) );
  CFD1XL \memory_reg[25][1]  ( .D(n649), .CP(clock), .Q(\memory[25][1] ), .QN(
        n121) );
  CFD1XL \memory_reg[25][0]  ( .D(n650), .CP(clock), .Q(\memory[25][0] ), .QN(
        n124) );
  CFD1XL \memory_reg[24][3]  ( .D(n651), .CP(clock), .Q(\memory[24][3] ), .QN(
        n129) );
  CFD1XL \memory_reg[24][2]  ( .D(n652), .CP(clock), .Q(\memory[24][2] ), .QN(
        n134) );
  CFD1XL \memory_reg[24][1]  ( .D(n653), .CP(clock), .Q(\memory[24][1] ), .QN(
        n137) );
  CFD1XL \memory_reg[24][0]  ( .D(n654), .CP(clock), .Q(\memory[24][0] ), .QN(
        n140) );
  CFD1XL \memory_reg[23][3]  ( .D(n655), .CP(clock), .Q(\memory[23][3] ), .QN(
        n145) );
  CFD1XL \memory_reg[23][2]  ( .D(n656), .CP(clock), .Q(\memory[23][2] ), .QN(
        n150) );
  CFD1XL \memory_reg[23][1]  ( .D(n657), .CP(clock), .Q(\memory[23][1] ), .QN(
        n153) );
  CFD1XL \memory_reg[23][0]  ( .D(n658), .CP(clock), .Q(\memory[23][0] ), .QN(
        n156) );
  CFD1XL \memory_reg[22][3]  ( .D(n659), .CP(clock), .Q(\memory[22][3] ), .QN(
        n162) );
  CFD1XL \memory_reg[22][2]  ( .D(n660), .CP(clock), .Q(\memory[22][2] ), .QN(
        n167) );
  CFD1XL \memory_reg[22][1]  ( .D(n661), .CP(clock), .Q(\memory[22][1] ), .QN(
        n170) );
  CFD1XL \memory_reg[22][0]  ( .D(n662), .CP(clock), .Q(\memory[22][0] ), .QN(
        n173) );
  CFD1XL \memory_reg[21][3]  ( .D(n663), .CP(clock), .Q(\memory[21][3] ), .QN(
        n177) );
  CFD1XL \memory_reg[21][2]  ( .D(n664), .CP(clock), .Q(\memory[21][2] ), .QN(
        n182) );
  CFD1XL \memory_reg[21][1]  ( .D(n665), .CP(clock), .Q(\memory[21][1] ), .QN(
        n185) );
  CFD1XL \memory_reg[21][0]  ( .D(n666), .CP(clock), .Q(\memory[21][0] ), .QN(
        n188) );
  CFD1XL \memory_reg[20][3]  ( .D(n667), .CP(clock), .Q(\memory[20][3] ), .QN(
        n192) );
  CFD1XL \memory_reg[20][2]  ( .D(n668), .CP(clock), .Q(\memory[20][2] ), .QN(
        n197) );
  CFD1XL \memory_reg[20][1]  ( .D(n669), .CP(clock), .Q(\memory[20][1] ), .QN(
        n200) );
  CFD1XL \memory_reg[20][0]  ( .D(n670), .CP(clock), .Q(\memory[20][0] ), .QN(
        n203) );
  CFD1XL \memory_reg[19][3]  ( .D(n671), .CP(clock), .Q(\memory[19][3] ), .QN(
        n207) );
  CFD1XL \memory_reg[19][2]  ( .D(n672), .CP(clock), .Q(\memory[19][2] ), .QN(
        n212) );
  CFD1XL \memory_reg[19][1]  ( .D(n673), .CP(clock), .Q(\memory[19][1] ), .QN(
        n215) );
  CFD1XL \memory_reg[19][0]  ( .D(n674), .CP(clock), .Q(\memory[19][0] ), .QN(
        n218) );
  CFD1XL \memory_reg[18][3]  ( .D(n675), .CP(clock), .Q(\memory[18][3] ), .QN(
        n222) );
  CFD1XL \memory_reg[18][2]  ( .D(n676), .CP(clock), .Q(\memory[18][2] ), .QN(
        n227) );
  CFD1XL \memory_reg[18][1]  ( .D(n677), .CP(clock), .Q(\memory[18][1] ), .QN(
        n230) );
  CFD1XL \memory_reg[18][0]  ( .D(n678), .CP(clock), .Q(\memory[18][0] ), .QN(
        n233) );
  CFD1XL \memory_reg[17][3]  ( .D(n679), .CP(clock), .Q(\memory[17][3] ), .QN(
        n237) );
  CFD1XL \memory_reg[17][2]  ( .D(n680), .CP(clock), .Q(\memory[17][2] ), .QN(
        n242) );
  CFD1XL \memory_reg[17][1]  ( .D(n681), .CP(clock), .Q(\memory[17][1] ), .QN(
        n245) );
  CFD1XL \memory_reg[17][0]  ( .D(n682), .CP(clock), .Q(\memory[17][0] ), .QN(
        n248) );
  CFD1XL \memory_reg[16][3]  ( .D(n683), .CP(clock), .Q(\memory[16][3] ), .QN(
        n252) );
  CFD1XL \memory_reg[16][2]  ( .D(n684), .CP(clock), .Q(\memory[16][2] ), .QN(
        n257) );
  CFD1XL \memory_reg[16][1]  ( .D(n685), .CP(clock), .Q(\memory[16][1] ), .QN(
        n260) );
  CFD1XL \memory_reg[16][0]  ( .D(n686), .CP(clock), .Q(\memory[16][0] ), .QN(
        n263) );
  CFD1XL \memory_reg[15][3]  ( .D(n687), .CP(clock), .Q(\memory[15][3] ), .QN(
        n268) );
  CFD1XL \memory_reg[15][2]  ( .D(n688), .CP(clock), .Q(\memory[15][2] ), .QN(
        n273) );
  CFD1XL \memory_reg[15][1]  ( .D(n689), .CP(clock), .Q(\memory[15][1] ), .QN(
        n276) );
  CFD1XL \memory_reg[15][0]  ( .D(n690), .CP(clock), .Q(\memory[15][0] ), .QN(
        n279) );
  CFD1XL \memory_reg[14][3]  ( .D(n691), .CP(clock), .Q(\memory[14][3] ), .QN(
        n284) );
  CFD1XL \memory_reg[14][2]  ( .D(n692), .CP(clock), .Q(\memory[14][2] ), .QN(
        n289) );
  CFD1XL \memory_reg[14][1]  ( .D(n693), .CP(clock), .Q(\memory[14][1] ), .QN(
        n292) );
  CFD1XL \memory_reg[14][0]  ( .D(n694), .CP(clock), .Q(\memory[14][0] ), .QN(
        n295) );
  CFD1XL \memory_reg[13][3]  ( .D(n695), .CP(clock), .Q(\memory[13][3] ), .QN(
        n299) );
  CFD1XL \memory_reg[13][2]  ( .D(n696), .CP(clock), .Q(\memory[13][2] ), .QN(
        n304) );
  CFD1XL \memory_reg[13][1]  ( .D(n697), .CP(clock), .Q(\memory[13][1] ), .QN(
        n307) );
  CFD1XL \memory_reg[13][0]  ( .D(n698), .CP(clock), .Q(\memory[13][0] ), .QN(
        n310) );
  CFD1XL \memory_reg[12][3]  ( .D(n699), .CP(clock), .Q(\memory[12][3] ), .QN(
        n314) );
  CFD1XL \memory_reg[12][2]  ( .D(n700), .CP(clock), .Q(\memory[12][2] ), .QN(
        n319) );
  CFD1XL \memory_reg[12][1]  ( .D(n701), .CP(clock), .Q(\memory[12][1] ), .QN(
        n322) );
  CFD1XL \memory_reg[12][0]  ( .D(n702), .CP(clock), .Q(\memory[12][0] ), .QN(
        n325) );
  CFD1XL \memory_reg[11][3]  ( .D(n703), .CP(clock), .Q(\memory[11][3] ), .QN(
        n329) );
  CFD1XL \memory_reg[11][2]  ( .D(n704), .CP(clock), .Q(\memory[11][2] ), .QN(
        n334) );
  CFD1XL \memory_reg[11][1]  ( .D(n705), .CP(clock), .Q(\memory[11][1] ), .QN(
        n337) );
  CFD1XL \memory_reg[11][0]  ( .D(n706), .CP(clock), .Q(\memory[11][0] ), .QN(
        n340) );
  CFD1XL \memory_reg[10][3]  ( .D(n707), .CP(clock), .Q(\memory[10][3] ), .QN(
        n344) );
  CFD1XL \memory_reg[10][2]  ( .D(n708), .CP(clock), .Q(\memory[10][2] ), .QN(
        n349) );
  CFD1XL \memory_reg[10][1]  ( .D(n709), .CP(clock), .Q(\memory[10][1] ), .QN(
        n352) );
  CFD1XL \memory_reg[10][0]  ( .D(n710), .CP(clock), .Q(\memory[10][0] ), .QN(
        n355) );
  CFD1XL \memory_reg[9][3]  ( .D(n711), .CP(clock), .Q(\memory[9][3] ), .QN(
        n359) );
  CFD1XL \memory_reg[9][2]  ( .D(n712), .CP(clock), .Q(\memory[9][2] ), .QN(
        n364) );
  CFD1XL \memory_reg[9][1]  ( .D(n713), .CP(clock), .Q(\memory[9][1] ), .QN(
        n367) );
  CFD1XL \memory_reg[9][0]  ( .D(n714), .CP(clock), .Q(\memory[9][0] ), .QN(
        n370) );
  CFD1XL \memory_reg[8][3]  ( .D(n715), .CP(clock), .Q(\memory[8][3] ), .QN(
        n374) );
  CFD1XL \memory_reg[8][2]  ( .D(n716), .CP(clock), .Q(\memory[8][2] ), .QN(
        n379) );
  CFD1XL \memory_reg[8][1]  ( .D(n717), .CP(clock), .Q(\memory[8][1] ), .QN(
        n382) );
  CFD1XL \memory_reg[8][0]  ( .D(n718), .CP(clock), .Q(\memory[8][0] ), .QN(
        n385) );
  CFD1XL \memory_reg[6][3]  ( .D(n723), .CP(clock), .Q(\memory[6][3] ), .QN(
        n406) );
  CFD1XL \memory_reg[6][2]  ( .D(n724), .CP(clock), .Q(\memory[6][2] ), .QN(
        n411) );
  CFD1XL \memory_reg[6][1]  ( .D(n725), .CP(clock), .Q(\memory[6][1] ), .QN(
        n414) );
  CFD1XL \memory_reg[6][0]  ( .D(n726), .CP(clock), .Q(\memory[6][0] ), .QN(
        n417) );
  CFD1XL \memory_reg[7][3]  ( .D(n719), .CP(clock), .Q(\memory[7][3] ), .QN(
        n390) );
  CFD1XL \memory_reg[7][2]  ( .D(n720), .CP(clock), .Q(\memory[7][2] ), .QN(
        n395) );
  CFD1XL \memory_reg[7][1]  ( .D(n721), .CP(clock), .Q(\memory[7][1] ), .QN(
        n398) );
  CFD1XL \memory_reg[7][0]  ( .D(n722), .CP(clock), .Q(\memory[7][0] ), .QN(
        n401) );
  CFD1XL \memory_reg[5][3]  ( .D(n727), .CP(clock), .Q(\memory[5][3] ), .QN(
        n423) );
  CFD1XL \memory_reg[5][2]  ( .D(n728), .CP(clock), .Q(\memory[5][2] ), .QN(
        n428) );
  CFD1XL \memory_reg[5][1]  ( .D(n729), .CP(clock), .Q(\memory[5][1] ), .QN(
        n431) );
  CFD1XL \memory_reg[5][0]  ( .D(n730), .CP(clock), .Q(\memory[5][0] ), .QN(
        n434) );
  CFD1XL \memory_reg[4][3]  ( .D(n731), .CP(clock), .Q(\memory[4][3] ), .QN(
        n439) );
  CFD1XL \memory_reg[4][2]  ( .D(n732), .CP(clock), .Q(\memory[4][2] ), .QN(
        n444) );
  CFD1XL \memory_reg[4][1]  ( .D(n733), .CP(clock), .Q(\memory[4][1] ), .QN(
        n447) );
  CFD1XL \memory_reg[4][0]  ( .D(n734), .CP(clock), .Q(\memory[4][0] ), .QN(
        n450) );
  CFD1XL \memory_reg[3][3]  ( .D(n735), .CP(clock), .Q(\memory[3][3] ), .QN(
        n454) );
  CFD1XL \memory_reg[3][2]  ( .D(n736), .CP(clock), .Q(\memory[3][2] ), .QN(
        n459) );
  CFD1XL \memory_reg[3][1]  ( .D(n737), .CP(clock), .Q(\memory[3][1] ), .QN(
        n462) );
  CFD1XL \memory_reg[2][3]  ( .D(n739), .CP(clock), .Q(\memory[2][3] ), .QN(
        n469) );
  CFD1XL \memory_reg[2][2]  ( .D(n740), .CP(clock), .Q(\memory[2][2] ), .QN(
        n474) );
  CFD1XL \memory_reg[2][1]  ( .D(n741), .CP(clock), .Q(\memory[2][1] ), .QN(
        n477) );
  CFD1XL \memory_reg[2][0]  ( .D(n742), .CP(clock), .Q(\memory[2][0] ), .QN(
        n480) );
  CFD1XL \memory_reg[3][0]  ( .D(n738), .CP(clock), .Q(\memory[3][0] ), .QN(
        n465) );
  CAOR2X4 U4 ( .A(empty), .B(n19), .C(n20), .D(n21), .Z(n626) );
  CND2XL U5 ( .A(n515), .B(reset), .Z(n498) );
  CANR2XL U6 ( .A(n527), .B(N121), .C(counter[30]), .D(n528), .Z(n526) );
  CDLY1XL U8 ( .A(counter[0]), .Z(n14) );
  COND3XL U9 ( .A(n533), .B(n524), .C(n534), .D(n535), .Z(n761) );
  COND3XL U356 ( .A(n523), .B(n524), .C(n525), .D(n526), .Z(n759) );
  COND1X1 U359 ( .A(n468), .B(n480), .C(n481), .Z(n742) );
  CIVX1 U362 ( .A(n504), .Z(n15) );
  CIVX2 U365 ( .A(n15), .Z(n791) );
  CIVX1 U387 ( .A(n47), .Z(n792) );
  CIVX2 U390 ( .A(n792), .Z(n793) );
  CIVX1 U393 ( .A(n68), .Z(n794) );
  CIVX2 U396 ( .A(n794), .Z(n795) );
  CIVX1 U403 ( .A(n84), .Z(n796) );
  CIVX2 U406 ( .A(n796), .Z(n797) );
  CIVX1 U409 ( .A(n100), .Z(n798) );
  CIVX2 U412 ( .A(n798), .Z(n799) );
  CIVX1 U419 ( .A(n116), .Z(n800) );
  CIVX2 U422 ( .A(n800), .Z(n801) );
  CIVX1 U425 ( .A(n132), .Z(n802) );
  CIVX2 U428 ( .A(n802), .Z(n803) );
  CIVX1 U435 ( .A(n148), .Z(n804) );
  CIVX2 U438 ( .A(n804), .Z(n805) );
  CIVX1 U441 ( .A(n165), .Z(n806) );
  CIVX2 U444 ( .A(n806), .Z(n807) );
  CIVX1 U451 ( .A(n180), .Z(n808) );
  CIVX2 U454 ( .A(n808), .Z(n809) );
  CIVX1 U457 ( .A(n195), .Z(n810) );
  CIVX2 U460 ( .A(n810), .Z(n811) );
  CIVX1 U461 ( .A(n210), .Z(n812) );
  CIVX2 U473 ( .A(n812), .Z(n813) );
  CIVX1 U480 ( .A(n225), .Z(n814) );
  CIVX2 U487 ( .A(n814), .Z(n815) );
  CIVX1 U497 ( .A(n240), .Z(n816) );
  CIVX2 U498 ( .A(n816), .Z(n817) );
  CIVX1 U502 ( .A(n255), .Z(n818) );
  CIVX2 U504 ( .A(n818), .Z(n819) );
  CIVX1 U516 ( .A(n271), .Z(n820) );
  CIVX2 U519 ( .A(n820), .Z(n821) );
  COND1X1 U520 ( .A(n389), .B(n390), .C(n391), .Z(n719) );
  COND1X1 U525 ( .A(n389), .B(n395), .C(n396), .Z(n720) );
  COND1X1 U609 ( .A(n389), .B(n398), .C(n399), .Z(n721) );
  CIVX1 U610 ( .A(n287), .Z(n822) );
  CIVX2 U614 ( .A(n822), .Z(n823) );
  CIVX1 U616 ( .A(n302), .Z(n824) );
  CIVX2 U618 ( .A(n824), .Z(n825) );
  CIVX1 U620 ( .A(n317), .Z(n826) );
  CIVX2 U621 ( .A(n826), .Z(n827) );
  CIVX1 U685 ( .A(n332), .Z(n828) );
  CIVX2 U686 ( .A(n828), .Z(n829) );
  CIVX1 U688 ( .A(n347), .Z(n830) );
  CIVX2 U696 ( .A(n830), .Z(n831) );
  CIVX1 U697 ( .A(n362), .Z(n832) );
  CIVX2 U698 ( .A(n832), .Z(n833) );
  CIVX1 U699 ( .A(n377), .Z(n834) );
  CIVX2 U700 ( .A(n834), .Z(n835) );
  COND1X1 U701 ( .A(n389), .B(n401), .C(n402), .Z(n722) );
  COND1X1 U702 ( .A(n422), .B(n423), .C(n424), .Z(n727) );
  COND1X1 U703 ( .A(n438), .B(n439), .C(n440), .Z(n731) );
  COND1X1 U704 ( .A(n453), .B(n454), .C(n455), .Z(n735) );
  COND1X1 U705 ( .A(n468), .B(n469), .C(n470), .Z(n739) );
  COND1X1 U706 ( .A(n483), .B(n484), .C(n485), .Z(n743) );
  COND1X1 U707 ( .A(n422), .B(n428), .C(n429), .Z(n728) );
  COND1X1 U708 ( .A(n438), .B(n444), .C(n445), .Z(n732) );
  COND1X1 U709 ( .A(n453), .B(n459), .C(n460), .Z(n736) );
  COND1X1 U710 ( .A(n468), .B(n474), .C(n475), .Z(n740) );
  COND1X1 U711 ( .A(n483), .B(n489), .C(n490), .Z(n744) );
  COND1X1 U712 ( .A(n422), .B(n431), .C(n432), .Z(n729) );
  COND1X1 U713 ( .A(n438), .B(n447), .C(n448), .Z(n733) );
  COND1X1 U714 ( .A(n453), .B(n462), .C(n463), .Z(n737) );
  COND1X1 U715 ( .A(n468), .B(n477), .C(n478), .Z(n741) );
  COND1X1 U716 ( .A(n483), .B(n492), .C(n493), .Z(n745) );
  CIVX1 U717 ( .A(n409), .Z(n836) );
  CIVX2 U718 ( .A(n836), .Z(n837) );
  COND1X1 U719 ( .A(n422), .B(n434), .C(n435), .Z(n730) );
  COND1X1 U720 ( .A(n438), .B(n450), .C(n451), .Z(n734) );
  COND1X1 U721 ( .A(n453), .B(n465), .C(n466), .Z(n738) );
  COND1X1 U722 ( .A(n483), .B(n495), .C(n496), .Z(n746) );
  CANR2XL U723 ( .A(N123), .B(n527), .C(counter[31]), .D(n528), .Z(n615) );
  CIVX2 U724 ( .A(n613), .Z(N248) );
  CANR2X2 U725 ( .A(N123), .B(n22), .C(n620), .D(counter[31]), .Z(n613) );
  COND4CX1 U726 ( .A(\memory[3][0] ), .B(n45), .C(n497), .D(n483), .Z(n496) );
  CIVXL U727 ( .A(rd_enable), .Z(n518) );
  COND3XL U728 ( .A(n613), .B(n524), .C(n614), .D(n615), .Z(n789) );
  CIVDXL U729 ( .A(N282), .Z0(n521) );
  COND1X1 U730 ( .A(n517), .B(n516), .C(rd_enable), .Z(n22) );
  CAOR1X2 U731 ( .A(n852), .B(n851), .C(N248), .Z(N282) );
  CNR2IX4 U732 ( .B(n17), .A(n528), .Z(n527) );
  CAN2X4 U733 ( .A(n17), .B(n515), .Z(n45) );
  CNR2X2 U734 ( .A(n619), .B(N282), .Z(n17) );
  CIVX4 U735 ( .A(n618), .Z(n528) );
  CANR1X1 U736 ( .A(n17), .B(n620), .C(N1652), .Z(n618) );
  CNR2X4 U737 ( .A(n528), .B(n21), .Z(n529) );
  COR6X1 U738 ( .A(counter[29]), .B(counter[28]), .C(counter[27]), .D(
        counter[9]), .E(counter[8]), .F(counter[30]), .Z(n847) );
  COR3X1 U739 ( .A(counter[14]), .B(counter[13]), .C(counter[12]), .Z(n845) );
  CANR3X1 U740 ( .A(counter[5]), .B(counter[4]), .C(counter[7]), .D(counter[6]), .Z(n843) );
  CIVX1 U741 ( .A(counter[5]), .Z(n842) );
  CIVX1 U742 ( .A(n843), .Z(n839) );
  CNR5X1 U743 ( .A(n14), .B(n839), .C(counter[1]), .D(counter[3]), .E(
        counter[2]), .Z(n841) );
  CNR2X1 U744 ( .A(counter[11]), .B(counter[10]), .Z(n840) );
  COND4CX1 U745 ( .A(n843), .B(n842), .C(n841), .D(n840), .Z(n844) );
  COR8X1 U746 ( .A(counter[17]), .B(counter[16]), .C(counter[15]), .D(
        counter[20]), .E(counter[19]), .F(counter[18]), .G(n845), .H(n844), 
        .Z(n846) );
  COR8X1 U747 ( .A(counter[23]), .B(counter[22]), .C(counter[21]), .D(
        counter[26]), .E(counter[25]), .F(counter[24]), .G(n847), .H(n846), 
        .Z(n848) );
  CND2IX1 U748 ( .B(counter[31]), .A(n848), .Z(N50) );
  COR6X1 U749 ( .A(N267), .B(N268), .C(N269), .D(N264), .E(N265), .F(N266), 
        .Z(n849) );
  CNR8X1 U750 ( .A(n849), .B(N263), .C(N261), .D(N262), .E(N257), .F(N258), 
        .G(N259), .H(N260), .Z(n852) );
  COR6X1 U751 ( .A(N254), .B(N255), .C(N256), .D(N251), .E(N252), .F(N253), 
        .Z(n850) );
  CNR8X1 U752 ( .A(n850), .B(N250), .C(N274), .D(N249), .E(N270), .F(N271), 
        .G(N272), .H(N273), .Z(n851) );
  fifo_DW01_sub_0 sub_42_aco ( .A(counter), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, rd_enable}), .CI(1'b0), .DIFF({N123, N121, N119, N117, 
        N115, N113, N111, N109, N107, N105, N103, N101, N99, N97, N95, N93, 
        N91, N89, N87, N85, N83, N81, N79, N77, N75, N73, N71, N69, N67, N65, 
        N63, N61}) );
  fifo_DW01_inc_0 add_74 ( .A({N248, N249, N250, N251, N252, N253, N254, N255, 
        N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
        N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279}), .SUM({N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, 
        N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, 
        N571, N570, N569, N568, N567, N566, N565, N564, N563}) );
  CFD1QXL \code_reg[3]  ( .D(n747), .CP(clock), .Q(code[3]) );
  CFD1QXL \code_reg[2]  ( .D(n749), .CP(clock), .Q(code[2]) );
  CFD1QXL \code_reg[1]  ( .D(n751), .CP(clock), .Q(code[1]) );
  CFD1QXL \code_reg[0]  ( .D(n753), .CP(clock), .Q(code[0]) );
  CFD1QXL \memory_reg[31][3]  ( .D(n755), .CP(clock), .Q(\memory[31][3] ) );
  CFD1QXL \memory_reg[31][2]  ( .D(n756), .CP(clock), .Q(\memory[31][2] ) );
  CFD1QXL \memory_reg[31][1]  ( .D(n757), .CP(clock), .Q(\memory[31][1] ) );
  CFD1QXL \memory_reg[31][0]  ( .D(n758), .CP(clock), .Q(\memory[31][0] ) );
endmodule


module decoder ( code, rd_enable, clock, BCD );
  input [3:0] code;
  output [7:0] BCD;
  input rd_enable, clock;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  assign BCD[7] = 1'b0;
  assign BCD[6] = 1'b0;
  assign BCD[5] = 1'b0;

  COND2X1 U4 ( .A(code[3]), .B(n3), .C(n4), .D(n5), .Z(n2) );
  COND11X1 U5 ( .A(n5), .B(n6), .C(n1), .D(n7), .Z(n13) );
  CND2X1 U6 ( .A(BCD[2]), .B(n1), .Z(n7) );
  CIVX1 U7 ( .A(n4), .Z(n6) );
  CIVX1 U8 ( .A(code[2]), .Z(n5) );
  COND11X1 U9 ( .A(n4), .B(code[2]), .C(n1), .D(n8), .Z(n14) );
  CND2X1 U10 ( .A(BCD[3]), .B(n1), .Z(n8) );
  CND2X1 U12 ( .A(code[3]), .B(n3), .Z(n4) );
  CIVX1 U13 ( .A(code[1]), .Z(n3) );
  COND1XL U14 ( .A(n9), .B(rd_enable), .C(n10), .Z(n15) );
  CFD1XL \BCD_reg[4]  ( .D(n15), .CP(clock), .Q(BCD[4]), .QN(n9) );
  CIVXL U2 ( .A(rd_enable), .Z(n1) );
  CAOR2XL U3 ( .A(BCD[1]), .B(n1), .C(rd_enable), .D(n2), .Z(n12) );
  COND3XL U11 ( .A(code[2]), .B(code[1]), .C(code[3]), .D(rd_enable), .Z(n10)
         );
  CAOR2XL U15 ( .A(rd_enable), .B(code[0]), .C(BCD[0]), .D(n1), .Z(n11) );
  CFD1QXL \BCD_reg[0]  ( .D(n11), .CP(clock), .Q(BCD[0]) );
  CFD1QXL \BCD_reg[3]  ( .D(n14), .CP(clock), .Q(BCD[3]) );
  CFD1QXL \BCD_reg[2]  ( .D(n13), .CP(clock), .Q(BCD[2]) );
  CFD1QXL \BCD_reg[1]  ( .D(n12), .CP(clock), .Q(BCD[1]) );
endmodule


module KSE ( clock, reset, row, read, BCD, valid, col );
  input [3:0] row;
  output [7:0] BCD;
  output [3:0] col;
  input clock, reset, read;
  output valid;
  wire   v, full, empty, wr_enable, rd_enable, n1, n2, n3, n4, n5, n6, n7;
  wire   [3:0] code;
  wire   [3:0] data;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;
  assign BCD[7] = 1'b0;
  assign BCD[6] = 1'b0;
  assign BCD[5] = 1'b0;

  CNIVXL U1 ( .A(read), .Z(n3) );
  CNIVX1 U2 ( .A(n2), .Z(n1) );
  CNIVX1 U3 ( .A(n3), .Z(n2) );
  CDLY1XL U4 ( .A(row[3]), .Z(n4) );
  CDLY1XL U5 ( .A(row[2]), .Z(n5) );
  CDLY1XL U6 ( .A(row[1]), .Z(n6) );
  CDLY1XL U7 ( .A(row[0]), .Z(n7) );
  keypad A ( .row({n4, n5, n6, n7}), .col(col), .data(data), .v(v), .clock(
        clock), .reset(reset) );
  controller B ( .v(v), .clock(clock), .reset(reset), .full(full), .empty(
        empty), .read(n1), .valid(valid), .wr_enable(wr_enable), .rd_enable(
        rd_enable) );
  fifo C ( .code(code), .full(full), .empty(empty), .data(data), .rd_enable(
        rd_enable), .wr_enable(wr_enable), .reset(reset), .clock(clock) );
  decoder D ( .code(code), .rd_enable(rd_enable), .clock(clock), .BCD({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, BCD[4:0]}) );
endmodule

